`timescale 1ns / 1ps


module 
 FIFO_36_2_166 #(parameter
///////////advanced parameters//////////
	DATA_WIDTH 					= 32,
	ADDRESS_BITS 				= 17,
///////////architecture parameters//////
	IFM_SIZE 					= 32,
	IFM_DEPTH 					= 3,
	KERNAL_SIZE 				= 6,
	NUMBER_OF_FILTERS 			= 6,
///////////generated parameters/////////
	IFM_SIZE_NEXT           	= IFM_SIZE - KERNAL_SIZE + 1,
	ADDRESS_SIZE_IFM        	= $clog2(IFM_SIZE*IFM_SIZE),
	ADDRESS_SIZE_NEXT_IFM   	= $clog2(IFM_SIZE_NEXT*IFM_SIZE_NEXT),
	ADDRESS_SIZE_WM         	= $clog2(IFM_DEPTH*NUMBER_OF_FILTERS),
	NUMBER_OF_IFM           	= IFM_DEPTH,      
	FIFO_SIZE               	= (KERNAL_SIZE-1)*IFM_SIZE + KERNAL_SIZE,
	NUMBER_OF_IFM_NEXT      	= NUMBER_OF_FILTERS,
	NUMBER_OF_WM            	= KERNAL_SIZE*KERNAL_SIZE,                              
	NUMBER_OF_BITS_SEL_IFM_NEXT = $clog2(NUMBER_OF_IFM_NEXT)
	)(
	input clk,
	input reset,
	input fifo_enable,
	input [DATA_WIDTH-1:0] fifo_data_in,
	input [DATA_WIDTH-1:0] fifo_data_in_2,
	output [DATA_WIDTH-1:0] fifo_data_out_1,
	output [DATA_WIDTH-1:0] fifo_data_out_2,
	output [DATA_WIDTH-1:0] fifo_data_out_3,
	output [DATA_WIDTH-1:0] fifo_data_out_4,
	output [DATA_WIDTH-1:0] fifo_data_out_5,
	output [DATA_WIDTH-1:0] fifo_data_out_6,
	output [DATA_WIDTH-1:0] fifo_data_out_7,
	output [DATA_WIDTH-1:0] fifo_data_out_8,
	output [DATA_WIDTH-1:0] fifo_data_out_9,
	output [DATA_WIDTH-1:0] fifo_data_out_10,
	output [DATA_WIDTH-1:0] fifo_data_out_11,
	output [DATA_WIDTH-1:0] fifo_data_out_12,
	output [DATA_WIDTH-1:0] fifo_data_out_13,
	output [DATA_WIDTH-1:0] fifo_data_out_14,
	output [DATA_WIDTH-1:0] fifo_data_out_15,
	output [DATA_WIDTH-1:0] fifo_data_out_16,
	output [DATA_WIDTH-1:0] fifo_data_out_17,
	output [DATA_WIDTH-1:0] fifo_data_out_18,
	output [DATA_WIDTH-1:0] fifo_data_out_19,
	output [DATA_WIDTH-1:0] fifo_data_out_20,
	output [DATA_WIDTH-1:0] fifo_data_out_21,
	output [DATA_WIDTH-1:0] fifo_data_out_22,
	output [DATA_WIDTH-1:0] fifo_data_out_23,
	output [DATA_WIDTH-1:0] fifo_data_out_24,
	output [DATA_WIDTH-1:0] fifo_data_out_25,
	output [DATA_WIDTH-1:0] fifo_data_out_26,
	output [DATA_WIDTH-1:0] fifo_data_out_27,
	output [DATA_WIDTH-1:0] fifo_data_out_28,
	output [DATA_WIDTH-1:0] fifo_data_out_29,
	output [DATA_WIDTH-1:0] fifo_data_out_30,
	output [DATA_WIDTH-1:0] fifo_data_out_31,
	output [DATA_WIDTH-1:0] fifo_data_out_32,
	output [DATA_WIDTH-1:0] fifo_data_out_33,
	output [DATA_WIDTH-1:0] fifo_data_out_34,
	output [DATA_WIDTH-1:0] fifo_data_out_35,
	output [DATA_WIDTH-1:0] fifo_data_out_36
	);
	reg	[DATA_WIDTH-1:0] FIFO  [FIFO_SIZE-1:0] ;
	always @ (posedge clk or posedge reset)
    begin
        if(reset)
		begin
			FIFO[0] <= 0;
			FIFO[1] <= 0;
			FIFO[2] <= 0;
			FIFO[3] <= 0;
			FIFO[4] <= 0;
			FIFO[5] <= 0;
			FIFO[6] <= 0;
			FIFO[7] <= 0;
			FIFO[8] <= 0;
			FIFO[9] <= 0;
			FIFO[10] <= 0;
			FIFO[11] <= 0;
			FIFO[12] <= 0;
			FIFO[13] <= 0;
			FIFO[14] <= 0;
			FIFO[15] <= 0;
			FIFO[16] <= 0;
			FIFO[17] <= 0;
			FIFO[18] <= 0;
			FIFO[19] <= 0;
			FIFO[20] <= 0;
			FIFO[21] <= 0;
			FIFO[22] <= 0;
			FIFO[23] <= 0;
			FIFO[24] <= 0;
			FIFO[25] <= 0;
			FIFO[26] <= 0;
			FIFO[27] <= 0;
			FIFO[28] <= 0;
			FIFO[29] <= 0;
			FIFO[30] <= 0;
			FIFO[31] <= 0;
			FIFO[32] <= 0;
			FIFO[33] <= 0;
			FIFO[34] <= 0;
			FIFO[35] <= 0;
			FIFO[36] <= 0;
			FIFO[37] <= 0;
			FIFO[38] <= 0;
			FIFO[39] <= 0;
			FIFO[40] <= 0;
			FIFO[41] <= 0;
			FIFO[42] <= 0;
			FIFO[43] <= 0;
			FIFO[44] <= 0;
			FIFO[45] <= 0;
			FIFO[46] <= 0;
			FIFO[47] <= 0;
			FIFO[48] <= 0;
			FIFO[49] <= 0;
			FIFO[50] <= 0;
			FIFO[51] <= 0;
			FIFO[52] <= 0;
			FIFO[53] <= 0;
			FIFO[54] <= 0;
			FIFO[55] <= 0;
			FIFO[56] <= 0;
			FIFO[57] <= 0;
			FIFO[58] <= 0;
			FIFO[59] <= 0;
			FIFO[60] <= 0;
			FIFO[61] <= 0;
			FIFO[62] <= 0;
			FIFO[63] <= 0;
			FIFO[64] <= 0;
			FIFO[65] <= 0;
			FIFO[66] <= 0;
			FIFO[67] <= 0;
			FIFO[68] <= 0;
			FIFO[69] <= 0;
			FIFO[70] <= 0;
			FIFO[71] <= 0;
			FIFO[72] <= 0;
			FIFO[73] <= 0;
			FIFO[74] <= 0;
			FIFO[75] <= 0;
			FIFO[76] <= 0;
			FIFO[77] <= 0;
			FIFO[78] <= 0;
			FIFO[79] <= 0;
			FIFO[80] <= 0;
			FIFO[81] <= 0;
			FIFO[82] <= 0;
			FIFO[83] <= 0;
			FIFO[84] <= 0;
			FIFO[85] <= 0;
			FIFO[86] <= 0;
			FIFO[87] <= 0;
			FIFO[88] <= 0;
			FIFO[89] <= 0;
			FIFO[90] <= 0;
			FIFO[91] <= 0;
			FIFO[92] <= 0;
			FIFO[93] <= 0;
			FIFO[94] <= 0;
			FIFO[95] <= 0;
			FIFO[96] <= 0;
			FIFO[97] <= 0;
			FIFO[98] <= 0;
			FIFO[99] <= 0;
			FIFO[100] <= 0;
			FIFO[101] <= 0;
			FIFO[102] <= 0;
			FIFO[103] <= 0;
			FIFO[104] <= 0;
			FIFO[105] <= 0;
			FIFO[106] <= 0;
			FIFO[107] <= 0;
			FIFO[108] <= 0;
			FIFO[109] <= 0;
			FIFO[110] <= 0;
			FIFO[111] <= 0;
			FIFO[112] <= 0;
			FIFO[113] <= 0;
			FIFO[114] <= 0;
			FIFO[115] <= 0;
			FIFO[116] <= 0;
			FIFO[117] <= 0;
			FIFO[118] <= 0;
			FIFO[119] <= 0;
			FIFO[120] <= 0;
			FIFO[121] <= 0;
			FIFO[122] <= 0;
			FIFO[123] <= 0;
			FIFO[124] <= 0;
			FIFO[125] <= 0;
			FIFO[126] <= 0;
			FIFO[127] <= 0;
			FIFO[128] <= 0;
			FIFO[129] <= 0;
			FIFO[130] <= 0;
			FIFO[131] <= 0;
			FIFO[132] <= 0;
			FIFO[133] <= 0;
			FIFO[134] <= 0;
			FIFO[135] <= 0;
			FIFO[136] <= 0;
			FIFO[137] <= 0;
			FIFO[138] <= 0;
			FIFO[139] <= 0;
			FIFO[140] <= 0;
			FIFO[141] <= 0;
			FIFO[142] <= 0;
			FIFO[143] <= 0;
			FIFO[144] <= 0;
			FIFO[145] <= 0;
			FIFO[146] <= 0;
			FIFO[147] <= 0;
			FIFO[148] <= 0;
			FIFO[149] <= 0;
			FIFO[150] <= 0;
			FIFO[151] <= 0;
			FIFO[152] <= 0;
			FIFO[153] <= 0;
			FIFO[154] <= 0;
			FIFO[155] <= 0;
			FIFO[156] <= 0;
			FIFO[157] <= 0;
			FIFO[158] <= 0;
			FIFO[159] <= 0;
			FIFO[160] <= 0;
			FIFO[161] <= 0;
			FIFO[162] <= 0;
			FIFO[163] <= 0;
			FIFO[164] <= 0;
			FIFO[165] <= 0;
		end
		else if(fifo_enable)
		begin
			FIFO[0] <= fifo_data_in_2;
			FIFO[1] <= fifo_data_in;
			FIFO[2] <= FIFO[0];
			FIFO[3] <= FIFO[1];
			FIFO[4] <= FIFO[2];
			FIFO[5] <= FIFO[3];
			FIFO[6] <= FIFO[4];
			FIFO[7] <= FIFO[5];
			FIFO[8] <= FIFO[6];
			FIFO[9] <= FIFO[7];
			FIFO[10] <= FIFO[8];
			FIFO[11] <= FIFO[9];
			FIFO[12] <= FIFO[10];
			FIFO[13] <= FIFO[11];
			FIFO[14] <= FIFO[12];
			FIFO[15] <= FIFO[13];
			FIFO[16] <= FIFO[14];
			FIFO[17] <= FIFO[15];
			FIFO[18] <= FIFO[16];
			FIFO[19] <= FIFO[17];
			FIFO[20] <= FIFO[18];
			FIFO[21] <= FIFO[19];
			FIFO[22] <= FIFO[20];
			FIFO[23] <= FIFO[21];
			FIFO[24] <= FIFO[22];
			FIFO[25] <= FIFO[23];
			FIFO[26] <= FIFO[24];
			FIFO[27] <= FIFO[25];
			FIFO[28] <= FIFO[26];
			FIFO[29] <= FIFO[27];
			FIFO[30] <= FIFO[28];
			FIFO[31] <= FIFO[29];
			FIFO[32] <= FIFO[30];
			FIFO[33] <= FIFO[31];
			FIFO[34] <= FIFO[32];
			FIFO[35] <= FIFO[33];
			FIFO[36] <= FIFO[34];
			FIFO[37] <= FIFO[35];
			FIFO[38] <= FIFO[36];
			FIFO[39] <= FIFO[37];
			FIFO[40] <= FIFO[38];
			FIFO[41] <= FIFO[39];
			FIFO[42] <= FIFO[40];
			FIFO[43] <= FIFO[41];
			FIFO[44] <= FIFO[42];
			FIFO[45] <= FIFO[43];
			FIFO[46] <= FIFO[44];
			FIFO[47] <= FIFO[45];
			FIFO[48] <= FIFO[46];
			FIFO[49] <= FIFO[47];
			FIFO[50] <= FIFO[48];
			FIFO[51] <= FIFO[49];
			FIFO[52] <= FIFO[50];
			FIFO[53] <= FIFO[51];
			FIFO[54] <= FIFO[52];
			FIFO[55] <= FIFO[53];
			FIFO[56] <= FIFO[54];
			FIFO[57] <= FIFO[55];
			FIFO[58] <= FIFO[56];
			FIFO[59] <= FIFO[57];
			FIFO[60] <= FIFO[58];
			FIFO[61] <= FIFO[59];
			FIFO[62] <= FIFO[60];
			FIFO[63] <= FIFO[61];
			FIFO[64] <= FIFO[62];
			FIFO[65] <= FIFO[63];
			FIFO[66] <= FIFO[64];
			FIFO[67] <= FIFO[65];
			FIFO[68] <= FIFO[66];
			FIFO[69] <= FIFO[67];
			FIFO[70] <= FIFO[68];
			FIFO[71] <= FIFO[69];
			FIFO[72] <= FIFO[70];
			FIFO[73] <= FIFO[71];
			FIFO[74] <= FIFO[72];
			FIFO[75] <= FIFO[73];
			FIFO[76] <= FIFO[74];
			FIFO[77] <= FIFO[75];
			FIFO[78] <= FIFO[76];
			FIFO[79] <= FIFO[77];
			FIFO[80] <= FIFO[78];
			FIFO[81] <= FIFO[79];
			FIFO[82] <= FIFO[80];
			FIFO[83] <= FIFO[81];
			FIFO[84] <= FIFO[82];
			FIFO[85] <= FIFO[83];
			FIFO[86] <= FIFO[84];
			FIFO[87] <= FIFO[85];
			FIFO[88] <= FIFO[86];
			FIFO[89] <= FIFO[87];
			FIFO[90] <= FIFO[88];
			FIFO[91] <= FIFO[89];
			FIFO[92] <= FIFO[90];
			FIFO[93] <= FIFO[91];
			FIFO[94] <= FIFO[92];
			FIFO[95] <= FIFO[93];
			FIFO[96] <= FIFO[94];
			FIFO[97] <= FIFO[95];
			FIFO[98] <= FIFO[96];
			FIFO[99] <= FIFO[97];
			FIFO[100] <= FIFO[98];
			FIFO[101] <= FIFO[99];
			FIFO[102] <= FIFO[100];
			FIFO[103] <= FIFO[101];
			FIFO[104] <= FIFO[102];
			FIFO[105] <= FIFO[103];
			FIFO[106] <= FIFO[104];
			FIFO[107] <= FIFO[105];
			FIFO[108] <= FIFO[106];
			FIFO[109] <= FIFO[107];
			FIFO[110] <= FIFO[108];
			FIFO[111] <= FIFO[109];
			FIFO[112] <= FIFO[110];
			FIFO[113] <= FIFO[111];
			FIFO[114] <= FIFO[112];
			FIFO[115] <= FIFO[113];
			FIFO[116] <= FIFO[114];
			FIFO[117] <= FIFO[115];
			FIFO[118] <= FIFO[116];
			FIFO[119] <= FIFO[117];
			FIFO[120] <= FIFO[118];
			FIFO[121] <= FIFO[119];
			FIFO[122] <= FIFO[120];
			FIFO[123] <= FIFO[121];
			FIFO[124] <= FIFO[122];
			FIFO[125] <= FIFO[123];
			FIFO[126] <= FIFO[124];
			FIFO[127] <= FIFO[125];
			FIFO[128] <= FIFO[126];
			FIFO[129] <= FIFO[127];
			FIFO[130] <= FIFO[128];
			FIFO[131] <= FIFO[129];
			FIFO[132] <= FIFO[130];
			FIFO[133] <= FIFO[131];
			FIFO[134] <= FIFO[132];
			FIFO[135] <= FIFO[133];
			FIFO[136] <= FIFO[134];
			FIFO[137] <= FIFO[135];
			FIFO[138] <= FIFO[136];
			FIFO[139] <= FIFO[137];
			FIFO[140] <= FIFO[138];
			FIFO[141] <= FIFO[139];
			FIFO[142] <= FIFO[140];
			FIFO[143] <= FIFO[141];
			FIFO[144] <= FIFO[142];
			FIFO[145] <= FIFO[143];
			FIFO[146] <= FIFO[144];
			FIFO[147] <= FIFO[145];
			FIFO[148] <= FIFO[146];
			FIFO[149] <= FIFO[147];
			FIFO[150] <= FIFO[148];
			FIFO[151] <= FIFO[149];
			FIFO[152] <= FIFO[150];
			FIFO[153] <= FIFO[151];
			FIFO[154] <= FIFO[152];
			FIFO[155] <= FIFO[153];
			FIFO[156] <= FIFO[154];
			FIFO[157] <= FIFO[155];
			FIFO[158] <= FIFO[156];
			FIFO[159] <= FIFO[157];
			FIFO[160] <= FIFO[158];
			FIFO[161] <= FIFO[159];
			FIFO[162] <= FIFO[160];
			FIFO[163] <= FIFO[161];
			FIFO[164] <= FIFO[162];
			FIFO[165] <= FIFO[163];
		end
	end

	assign    fifo_data_out_1 = FIFO[(KERNAL_SIZE-1)*IFM_SIZE+(KERNAL_SIZE-1)];
	assign    fifo_data_out_2 = FIFO[(KERNAL_SIZE-1)*IFM_SIZE+(KERNAL_SIZE-2)];
	assign    fifo_data_out_3 = FIFO[(KERNAL_SIZE-1)*IFM_SIZE+(KERNAL_SIZE-3)];
	assign    fifo_data_out_4 = FIFO[(KERNAL_SIZE-1)*IFM_SIZE+(KERNAL_SIZE-4)];
	assign    fifo_data_out_5 = FIFO[(KERNAL_SIZE-1)*IFM_SIZE+(KERNAL_SIZE-5)];
	assign    fifo_data_out_6 = FIFO[(KERNAL_SIZE-1)*IFM_SIZE+(KERNAL_SIZE-6)];
	
	assign    fifo_data_out_7 = FIFO[(KERNAL_SIZE-2)*IFM_SIZE+(KERNAL_SIZE-1)];
	assign    fifo_data_out_8 = FIFO[(KERNAL_SIZE-2)*IFM_SIZE+(KERNAL_SIZE-2)];
	assign    fifo_data_out_9 = FIFO[(KERNAL_SIZE-2)*IFM_SIZE+(KERNAL_SIZE-3)];
	assign    fifo_data_out_10 = FIFO[(KERNAL_SIZE-2)*IFM_SIZE+(KERNAL_SIZE-4)];
	assign    fifo_data_out_11 = FIFO[(KERNAL_SIZE-2)*IFM_SIZE+(KERNAL_SIZE-5)];
	assign    fifo_data_out_12 = FIFO[(KERNAL_SIZE-2)*IFM_SIZE+(KERNAL_SIZE-6)];
	
	assign    fifo_data_out_13 = FIFO[(KERNAL_SIZE-3)*IFM_SIZE+(KERNAL_SIZE-1)];
	assign    fifo_data_out_14 = FIFO[(KERNAL_SIZE-3)*IFM_SIZE+(KERNAL_SIZE-2)];
	assign    fifo_data_out_15 = FIFO[(KERNAL_SIZE-3)*IFM_SIZE+(KERNAL_SIZE-3)];
	assign    fifo_data_out_16 = FIFO[(KERNAL_SIZE-3)*IFM_SIZE+(KERNAL_SIZE-4)];
	assign    fifo_data_out_17 = FIFO[(KERNAL_SIZE-3)*IFM_SIZE+(KERNAL_SIZE-5)];
	assign    fifo_data_out_18 = FIFO[(KERNAL_SIZE-3)*IFM_SIZE+(KERNAL_SIZE-6)];
	
	assign    fifo_data_out_19 = FIFO[(KERNAL_SIZE-4)*IFM_SIZE+(KERNAL_SIZE-1)];
	assign    fifo_data_out_20 = FIFO[(KERNAL_SIZE-4)*IFM_SIZE+(KERNAL_SIZE-2)];
	assign    fifo_data_out_21 = FIFO[(KERNAL_SIZE-4)*IFM_SIZE+(KERNAL_SIZE-3)];
	assign    fifo_data_out_22 = FIFO[(KERNAL_SIZE-4)*IFM_SIZE+(KERNAL_SIZE-4)];
	assign    fifo_data_out_23 = FIFO[(KERNAL_SIZE-4)*IFM_SIZE+(KERNAL_SIZE-5)];
	assign    fifo_data_out_24 = FIFO[(KERNAL_SIZE-4)*IFM_SIZE+(KERNAL_SIZE-6)];
	
	assign    fifo_data_out_25 = FIFO[(KERNAL_SIZE-5)*IFM_SIZE+(KERNAL_SIZE-1)];
	assign    fifo_data_out_26 = FIFO[(KERNAL_SIZE-5)*IFM_SIZE+(KERNAL_SIZE-2)];
	assign    fifo_data_out_27 = FIFO[(KERNAL_SIZE-5)*IFM_SIZE+(KERNAL_SIZE-3)];
	assign    fifo_data_out_28 = FIFO[(KERNAL_SIZE-5)*IFM_SIZE+(KERNAL_SIZE-4)];
	assign    fifo_data_out_29 = FIFO[(KERNAL_SIZE-5)*IFM_SIZE+(KERNAL_SIZE-5)];
	assign    fifo_data_out_30 = FIFO[(KERNAL_SIZE-5)*IFM_SIZE+(KERNAL_SIZE-6)];
	
	assign    fifo_data_out_31 = FIFO[(KERNAL_SIZE-6)*IFM_SIZE+(KERNAL_SIZE-1)];
	assign    fifo_data_out_32 = FIFO[(KERNAL_SIZE-6)*IFM_SIZE+(KERNAL_SIZE-2)];
	assign    fifo_data_out_33 = FIFO[(KERNAL_SIZE-6)*IFM_SIZE+(KERNAL_SIZE-3)];
	assign    fifo_data_out_34 = FIFO[(KERNAL_SIZE-6)*IFM_SIZE+(KERNAL_SIZE-4)];
	assign    fifo_data_out_35 = FIFO[(KERNAL_SIZE-6)*IFM_SIZE+(KERNAL_SIZE-5)];
	assign    fifo_data_out_36 = FIFO[(KERNAL_SIZE-6)*IFM_SIZE+(KERNAL_SIZE-6)];
	
endmodule