`timescale 1ns / 1ps


module 
 Float_Divider #(parameter
	DATA_WIDTH = 32
	,E = 8
	,M = 23
	)(
	input [DATA_WIDTH - 1:0] in1,
	input [DATA_WIDTH - 1:0] in2,
	output [DATA_WIDTH - 1:0] out
	);
	wire  [DATA_WIDTH - 1:0] in2_rec;
	 
	assign  in2_rec =   (in2 == 32'b 01000000100000000000000000000000) ? (32'b 00111110100000000000000000000000) :
						(in2 == 32'b 01000001000100000000000000000000) ? (32'b 00111101111000111000110110100100) :
						(in2 == 32'b 01000001100000000000000000000000) ? (32'b 00111101100000000000000000000000) :
						(in2 == 32'b 01000001110010000000000000000000) ? (32'b 00111101001000111101011100001010) :
						(32'b 00111100111000111011110011010011);
	
	Float_Multiplier #(.DATA_WIDTH(DATA_WIDTH), .E(E), .M(M))	M1 ( .in1 (in1) ,.in2 (in2_rec),.out(out));
	

endmodule
