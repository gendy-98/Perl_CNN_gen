`timescale 1ns / 1ps


module 
 top_fcA_1 #(parameter
///////////advanced parameters//////////
	DATA_WIDTH 					= 32,
///////////architecture parameters//////
	IFM_SIZE              = 1,
	IFM_DEPTH				= 160,
	//////////////////////////////////////
    ADDRESS_BITS        = 17,
    ARITH_TYPE          = 0,
    ADDRESS_SIZE_IFM        = $clog2(IFM_SIZE*IFM_SIZE),
    ADDRESS_SIZE_WM        = $clog2(IFM_DEPTH),
    NUMBER_OF_WM        = 100

	)(
	input clk,
	input reset,
    /////////////////////////////////////////////////////
    input [DATA_WIDTH-1:0]   riscv_data,
	input [ADDRESS_BITS-1:0] riscv_address,
	/////////////////////////////////////////////////////
	input [NUMBER_OF_WM-1:0] wm_enable_write,
	input  bm_enable_write,
    /////////////////////////////////////////////////////	 
    input [DATA_WIDTH-1:0] data_in_from_previous,	 
	input  start_from_previous,  
    output end_to_previous,
    output enable_read_current,
    output enable_write_next,

    output bias_sel,
    
    ////////////////////////////////////////// for next  
    output start_to_next,
    output [DATA_WIDTH-1:0]   reg_out_FC_1 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_2 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_3 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_4 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_5 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_6 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_7 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_8 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_9 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_10 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_11 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_12 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_13 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_14 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_15 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_16 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_17 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_18 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_19 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_20 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_21 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_22 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_23 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_24 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_25 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_26 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_27 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_28 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_29 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_30 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_31 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_32 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_33 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_34 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_35 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_36 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_37 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_38 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_39 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_40 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_41 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_42 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_43 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_44 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_45 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_46 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_47 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_48 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_49 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_50 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_51 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_52 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_53 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_54 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_55 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_56 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_57 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_58 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_59 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_60 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_61 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_62 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_63 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_64 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_65 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_66 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_67 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_68 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_69 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_70 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_71 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_72 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_73 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_74 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_75 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_76 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_77 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_78 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_79 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_80 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_81 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_82 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_83 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_84 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_85 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_86 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_87 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_88 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_89 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_90 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_91 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_92 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_93 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_94 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_95 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_96 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_97 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_98 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_99 ,
    output [DATA_WIDTH-1:0]   reg_out_FC_100 ,
    output [DATA_WIDTH-1:0]   data_bias_1 ,
    output [DATA_WIDTH-1:0]   data_bias_2 ,
    output [DATA_WIDTH-1:0]   data_bias_3 ,
    output [DATA_WIDTH-1:0]   data_bias_4 ,
    output [DATA_WIDTH-1:0]   data_bias_5 ,
    output [DATA_WIDTH-1:0]   data_bias_6 ,
    output [DATA_WIDTH-1:0]   data_bias_7 ,
    output [DATA_WIDTH-1:0]   data_bias_8 ,
    output [DATA_WIDTH-1:0]   data_bias_9 ,
    output [DATA_WIDTH-1:0]   data_bias_10 ,
    output [DATA_WIDTH-1:0]   data_bias_11 ,
    output [DATA_WIDTH-1:0]   data_bias_12 ,
    output [DATA_WIDTH-1:0]   data_bias_13 ,
    output [DATA_WIDTH-1:0]   data_bias_14 ,
    output [DATA_WIDTH-1:0]   data_bias_15 ,
    output [DATA_WIDTH-1:0]   data_bias_16 ,
    output [DATA_WIDTH-1:0]   data_bias_17 ,
    output [DATA_WIDTH-1:0]   data_bias_18 ,
    output [DATA_WIDTH-1:0]   data_bias_19 ,
    output [DATA_WIDTH-1:0]   data_bias_20 ,
    output [DATA_WIDTH-1:0]   data_bias_21 ,
    output [DATA_WIDTH-1:0]   data_bias_22 ,
    output [DATA_WIDTH-1:0]   data_bias_23 ,
    output [DATA_WIDTH-1:0]   data_bias_24 ,
    output [DATA_WIDTH-1:0]   data_bias_25 ,
    output [DATA_WIDTH-1:0]   data_bias_26 ,
    output [DATA_WIDTH-1:0]   data_bias_27 ,
    output [DATA_WIDTH-1:0]   data_bias_28 ,
    output [DATA_WIDTH-1:0]   data_bias_29 ,
    output [DATA_WIDTH-1:0]   data_bias_30 ,
    output [DATA_WIDTH-1:0]   data_bias_31 ,
    output [DATA_WIDTH-1:0]   data_bias_32 ,
    output [DATA_WIDTH-1:0]   data_bias_33 ,
    output [DATA_WIDTH-1:0]   data_bias_34 ,
    output [DATA_WIDTH-1:0]   data_bias_35 ,
    output [DATA_WIDTH-1:0]   data_bias_36 ,
    output [DATA_WIDTH-1:0]   data_bias_37 ,
    output [DATA_WIDTH-1:0]   data_bias_38 ,
    output [DATA_WIDTH-1:0]   data_bias_39 ,
    output [DATA_WIDTH-1:0]   data_bias_40 ,
    output [DATA_WIDTH-1:0]   data_bias_41 ,
    output [DATA_WIDTH-1:0]   data_bias_42 ,
    output [DATA_WIDTH-1:0]   data_bias_43 ,
    output [DATA_WIDTH-1:0]   data_bias_44 ,
    output [DATA_WIDTH-1:0]   data_bias_45 ,
    output [DATA_WIDTH-1:0]   data_bias_46 ,
    output [DATA_WIDTH-1:0]   data_bias_47 ,
    output [DATA_WIDTH-1:0]   data_bias_48 ,
    output [DATA_WIDTH-1:0]   data_bias_49 ,
    output [DATA_WIDTH-1:0]   data_bias_50 ,
    output [DATA_WIDTH-1:0]   data_bias_51 ,
    output [DATA_WIDTH-1:0]   data_bias_52 ,
    output [DATA_WIDTH-1:0]   data_bias_53 ,
    output [DATA_WIDTH-1:0]   data_bias_54 ,
    output [DATA_WIDTH-1:0]   data_bias_55 ,
    output [DATA_WIDTH-1:0]   data_bias_56 ,
    output [DATA_WIDTH-1:0]   data_bias_57 ,
    output [DATA_WIDTH-1:0]   data_bias_58 ,
    output [DATA_WIDTH-1:0]   data_bias_59 ,
    output [DATA_WIDTH-1:0]   data_bias_60 ,
    output [DATA_WIDTH-1:0]   data_bias_61 ,
    output [DATA_WIDTH-1:0]   data_bias_62 ,
    output [DATA_WIDTH-1:0]   data_bias_63 ,
    output [DATA_WIDTH-1:0]   data_bias_64 ,
    output [DATA_WIDTH-1:0]   data_bias_65 ,
    output [DATA_WIDTH-1:0]   data_bias_66 ,
    output [DATA_WIDTH-1:0]   data_bias_67 ,
    output [DATA_WIDTH-1:0]   data_bias_68 ,
    output [DATA_WIDTH-1:0]   data_bias_69 ,
    output [DATA_WIDTH-1:0]   data_bias_70 ,
    output [DATA_WIDTH-1:0]   data_bias_71 ,
    output [DATA_WIDTH-1:0]   data_bias_72 ,
    output [DATA_WIDTH-1:0]   data_bias_73 ,
    output [DATA_WIDTH-1:0]   data_bias_74 ,
    output [DATA_WIDTH-1:0]   data_bias_75 ,
    output [DATA_WIDTH-1:0]   data_bias_76 ,
    output [DATA_WIDTH-1:0]   data_bias_77 ,
    output [DATA_WIDTH-1:0]   data_bias_78 ,
    output [DATA_WIDTH-1:0]   data_bias_79 ,
    output [DATA_WIDTH-1:0]   data_bias_80 ,
    output [DATA_WIDTH-1:0]   data_bias_81 ,
    output [DATA_WIDTH-1:0]   data_bias_82 ,
    output [DATA_WIDTH-1:0]   data_bias_83 ,
    output [DATA_WIDTH-1:0]   data_bias_84 ,
    output [DATA_WIDTH-1:0]   data_bias_85 ,
    output [DATA_WIDTH-1:0]   data_bias_86 ,
    output [DATA_WIDTH-1:0]   data_bias_87 ,
    output [DATA_WIDTH-1:0]   data_bias_88 ,
    output [DATA_WIDTH-1:0]   data_bias_89 ,
    output [DATA_WIDTH-1:0]   data_bias_90 ,
    output [DATA_WIDTH-1:0]   data_bias_91 ,
    output [DATA_WIDTH-1:0]   data_bias_92 ,
    output [DATA_WIDTH-1:0]   data_bias_93 ,
    output [DATA_WIDTH-1:0]   data_bias_94 ,
    output [DATA_WIDTH-1:0]   data_bias_95 ,
    output [DATA_WIDTH-1:0]   data_bias_96 ,
    output [DATA_WIDTH-1:0]   data_bias_97 ,
    output [DATA_WIDTH-1:0]   data_bias_98 ,
    output [DATA_WIDTH-1:0]   data_bias_99 ,
    output [DATA_WIDTH-1:0]   data_bias_100 ,
	input  end_from_next
	);

    wire wm_enable_read;
    wire wm_addr_sel;
    wire [ADDRESS_SIZE_WM-1:0] wm_address_read_current;  
    
    wire fc_output_ready;


	FCA1_CU #(
    .IFM_DEPTH(IFM_DEPTH)) 
    CU
    (
    .clk(clk),
    .reset(reset),
	.start_from_previous(start_from_previous), 
	.end_from_next(end_from_next),
	.wm_addr_sel(wm_addr_sel),
    .wm_enable_read (wm_enable_read),
    .wm_address_read_current(wm_address_read_current), 
	.enable_read_current(enable_read_current),
    .end_to_previous (end_to_previous),    
    .enable_write_next (enable_write_next),
    .fc_output_ready (fc_output_ready),
    .bias_sel(bias_sel),
    .start_to_next (start_to_next)  
   );

	FCA1_DP #(.DATA_WIDTH(DATA_WIDTH), .ARITH_TYPE(ARITH_TYPE),
    .IFM_DEPTH(IFM_DEPTH), .NUMBER_OF_WM(NUMBER_OF_WM)) 
    DP
	(
    .clk(clk),
	.reset(reset),	
	.riscv_data(riscv_data),
	.riscv_address(riscv_address),
	/////////////////////////////////
    .wm_addr_sel (wm_addr_sel) , 
    .wm_enable_read (wm_enable_read),
    .wm_enable_write (wm_enable_write),
    .wm_address_read_current (wm_address_read_current),
    ///////////////////////////////////
    .bm_enable_write (bm_enable_write),
    ///////////////////////////////////
	.data_in_from_previous(data_in_from_previous),
	
	/////////////////////////////////////
   
    .reg_out_FC_1(reg_out_FC_1) , 
    .reg_out_FC_2(reg_out_FC_2) , 
    .reg_out_FC_3(reg_out_FC_3) , 
    .reg_out_FC_4(reg_out_FC_4) , 
    .reg_out_FC_5(reg_out_FC_5) , 
    .reg_out_FC_6(reg_out_FC_6) , 
    .reg_out_FC_7(reg_out_FC_7) , 
    .reg_out_FC_8(reg_out_FC_8) , 
    .reg_out_FC_9(reg_out_FC_9) , 
    .reg_out_FC_10(reg_out_FC_10) , 
    .reg_out_FC_11(reg_out_FC_11) , 
    .reg_out_FC_12(reg_out_FC_12) , 
    .reg_out_FC_13(reg_out_FC_13) , 
    .reg_out_FC_14(reg_out_FC_14) , 
    .reg_out_FC_15(reg_out_FC_15) , 
    .reg_out_FC_16(reg_out_FC_16) , 
    .reg_out_FC_17(reg_out_FC_17) , 
    .reg_out_FC_18(reg_out_FC_18) , 
    .reg_out_FC_19(reg_out_FC_19) , 
    .reg_out_FC_20(reg_out_FC_20) , 
    .reg_out_FC_21(reg_out_FC_21) , 
    .reg_out_FC_22(reg_out_FC_22) , 
    .reg_out_FC_23(reg_out_FC_23) , 
    .reg_out_FC_24(reg_out_FC_24) , 
    .reg_out_FC_25(reg_out_FC_25) , 
    .reg_out_FC_26(reg_out_FC_26) , 
    .reg_out_FC_27(reg_out_FC_27) , 
    .reg_out_FC_28(reg_out_FC_28) , 
    .reg_out_FC_29(reg_out_FC_29) , 
    .reg_out_FC_30(reg_out_FC_30) , 
    .reg_out_FC_31(reg_out_FC_31) , 
    .reg_out_FC_32(reg_out_FC_32) , 
    .reg_out_FC_33(reg_out_FC_33) , 
    .reg_out_FC_34(reg_out_FC_34) , 
    .reg_out_FC_35(reg_out_FC_35) , 
    .reg_out_FC_36(reg_out_FC_36) , 
    .reg_out_FC_37(reg_out_FC_37) , 
    .reg_out_FC_38(reg_out_FC_38) , 
    .reg_out_FC_39(reg_out_FC_39) , 
    .reg_out_FC_40(reg_out_FC_40) , 
    .reg_out_FC_41(reg_out_FC_41) , 
    .reg_out_FC_42(reg_out_FC_42) , 
    .reg_out_FC_43(reg_out_FC_43) , 
    .reg_out_FC_44(reg_out_FC_44) , 
    .reg_out_FC_45(reg_out_FC_45) , 
    .reg_out_FC_46(reg_out_FC_46) , 
    .reg_out_FC_47(reg_out_FC_47) , 
    .reg_out_FC_48(reg_out_FC_48) , 
    .reg_out_FC_49(reg_out_FC_49) , 
    .reg_out_FC_50(reg_out_FC_50) , 
    .reg_out_FC_51(reg_out_FC_51) , 
    .reg_out_FC_52(reg_out_FC_52) , 
    .reg_out_FC_53(reg_out_FC_53) , 
    .reg_out_FC_54(reg_out_FC_54) , 
    .reg_out_FC_55(reg_out_FC_55) , 
    .reg_out_FC_56(reg_out_FC_56) , 
    .reg_out_FC_57(reg_out_FC_57) , 
    .reg_out_FC_58(reg_out_FC_58) , 
    .reg_out_FC_59(reg_out_FC_59) , 
    .reg_out_FC_60(reg_out_FC_60) , 
    .reg_out_FC_61(reg_out_FC_61) , 
    .reg_out_FC_62(reg_out_FC_62) , 
    .reg_out_FC_63(reg_out_FC_63) , 
    .reg_out_FC_64(reg_out_FC_64) , 
    .reg_out_FC_65(reg_out_FC_65) , 
    .reg_out_FC_66(reg_out_FC_66) , 
    .reg_out_FC_67(reg_out_FC_67) , 
    .reg_out_FC_68(reg_out_FC_68) , 
    .reg_out_FC_69(reg_out_FC_69) , 
    .reg_out_FC_70(reg_out_FC_70) , 
    .reg_out_FC_71(reg_out_FC_71) , 
    .reg_out_FC_72(reg_out_FC_72) , 
    .reg_out_FC_73(reg_out_FC_73) , 
    .reg_out_FC_74(reg_out_FC_74) , 
    .reg_out_FC_75(reg_out_FC_75) , 
    .reg_out_FC_76(reg_out_FC_76) , 
    .reg_out_FC_77(reg_out_FC_77) , 
    .reg_out_FC_78(reg_out_FC_78) , 
    .reg_out_FC_79(reg_out_FC_79) , 
    .reg_out_FC_80(reg_out_FC_80) , 
    .reg_out_FC_81(reg_out_FC_81) , 
    .reg_out_FC_82(reg_out_FC_82) , 
    .reg_out_FC_83(reg_out_FC_83) , 
    .reg_out_FC_84(reg_out_FC_84) , 
    .reg_out_FC_85(reg_out_FC_85) , 
    .reg_out_FC_86(reg_out_FC_86) , 
    .reg_out_FC_87(reg_out_FC_87) , 
    .reg_out_FC_88(reg_out_FC_88) , 
    .reg_out_FC_89(reg_out_FC_89) , 
    .reg_out_FC_90(reg_out_FC_90) , 
    .reg_out_FC_91(reg_out_FC_91) , 
    .reg_out_FC_92(reg_out_FC_92) , 
    .reg_out_FC_93(reg_out_FC_93) , 
    .reg_out_FC_94(reg_out_FC_94) , 
    .reg_out_FC_95(reg_out_FC_95) , 
    .reg_out_FC_96(reg_out_FC_96) , 
    .reg_out_FC_97(reg_out_FC_97) , 
    .reg_out_FC_98(reg_out_FC_98) , 
    .reg_out_FC_99(reg_out_FC_99) , 
    .reg_out_FC_100(reg_out_FC_100) , 
    .data_bias_1  (data_bias_1 ),
    .data_bias_2  (data_bias_2 ),
    .data_bias_3  (data_bias_3 ),
    .data_bias_4  (data_bias_4 ),
    .data_bias_5  (data_bias_5 ),
    .data_bias_6  (data_bias_6 ),
    .data_bias_7  (data_bias_7 ),
    .data_bias_8  (data_bias_8 ),
    .data_bias_9  (data_bias_9 ),
    .data_bias_10  (data_bias_10 ),
    .data_bias_11  (data_bias_11 ),
    .data_bias_12  (data_bias_12 ),
    .data_bias_13  (data_bias_13 ),
    .data_bias_14  (data_bias_14 ),
    .data_bias_15  (data_bias_15 ),
    .data_bias_16  (data_bias_16 ),
    .data_bias_17  (data_bias_17 ),
    .data_bias_18  (data_bias_18 ),
    .data_bias_19  (data_bias_19 ),
    .data_bias_20  (data_bias_20 ),
    .data_bias_21  (data_bias_21 ),
    .data_bias_22  (data_bias_22 ),
    .data_bias_23  (data_bias_23 ),
    .data_bias_24  (data_bias_24 ),
    .data_bias_25  (data_bias_25 ),
    .data_bias_26  (data_bias_26 ),
    .data_bias_27  (data_bias_27 ),
    .data_bias_28  (data_bias_28 ),
    .data_bias_29  (data_bias_29 ),
    .data_bias_30  (data_bias_30 ),
    .data_bias_31  (data_bias_31 ),
    .data_bias_32  (data_bias_32 ),
    .data_bias_33  (data_bias_33 ),
    .data_bias_34  (data_bias_34 ),
    .data_bias_35  (data_bias_35 ),
    .data_bias_36  (data_bias_36 ),
    .data_bias_37  (data_bias_37 ),
    .data_bias_38  (data_bias_38 ),
    .data_bias_39  (data_bias_39 ),
    .data_bias_40  (data_bias_40 ),
    .data_bias_41  (data_bias_41 ),
    .data_bias_42  (data_bias_42 ),
    .data_bias_43  (data_bias_43 ),
    .data_bias_44  (data_bias_44 ),
    .data_bias_45  (data_bias_45 ),
    .data_bias_46  (data_bias_46 ),
    .data_bias_47  (data_bias_47 ),
    .data_bias_48  (data_bias_48 ),
    .data_bias_49  (data_bias_49 ),
    .data_bias_50  (data_bias_50 ),
    .data_bias_51  (data_bias_51 ),
    .data_bias_52  (data_bias_52 ),
    .data_bias_53  (data_bias_53 ),
    .data_bias_54  (data_bias_54 ),
    .data_bias_55  (data_bias_55 ),
    .data_bias_56  (data_bias_56 ),
    .data_bias_57  (data_bias_57 ),
    .data_bias_58  (data_bias_58 ),
    .data_bias_59  (data_bias_59 ),
    .data_bias_60  (data_bias_60 ),
    .data_bias_61  (data_bias_61 ),
    .data_bias_62  (data_bias_62 ),
    .data_bias_63  (data_bias_63 ),
    .data_bias_64  (data_bias_64 ),
    .data_bias_65  (data_bias_65 ),
    .data_bias_66  (data_bias_66 ),
    .data_bias_67  (data_bias_67 ),
    .data_bias_68  (data_bias_68 ),
    .data_bias_69  (data_bias_69 ),
    .data_bias_70  (data_bias_70 ),
    .data_bias_71  (data_bias_71 ),
    .data_bias_72  (data_bias_72 ),
    .data_bias_73  (data_bias_73 ),
    .data_bias_74  (data_bias_74 ),
    .data_bias_75  (data_bias_75 ),
    .data_bias_76  (data_bias_76 ),
    .data_bias_77  (data_bias_77 ),
    .data_bias_78  (data_bias_78 ),
    .data_bias_79  (data_bias_79 ),
    .data_bias_80  (data_bias_80 ),
    .data_bias_81  (data_bias_81 ),
    .data_bias_82  (data_bias_82 ),
    .data_bias_83  (data_bias_83 ),
    .data_bias_84  (data_bias_84 ),
    .data_bias_85  (data_bias_85 ),
    .data_bias_86  (data_bias_86 ),
    .data_bias_87  (data_bias_87 ),
    .data_bias_88  (data_bias_88 ),
    .data_bias_89  (data_bias_89 ),
    .data_bias_90  (data_bias_90 ),
    .data_bias_91  (data_bias_91 ),
    .data_bias_92  (data_bias_92 ),
    .data_bias_93  (data_bias_93 ),
    .data_bias_94  (data_bias_94 ),
    .data_bias_95  (data_bias_95 ),
    .data_bias_96  (data_bias_96 ),
    .data_bias_97  (data_bias_97 ),
    .data_bias_98  (data_bias_98 ),
    .data_bias_99  (data_bias_99 ),
    .data_bias_100  (data_bias_100 ),
    .fc_output_ready (fc_output_ready)
	);
endmodule
