`timescale 1ns / 1ps


module 
 Fixed_Divider #(parameter
	DATA_WIDTH = 32
	,E = 8
	,M = 27
	)(
	input [DATA_WIDTH - 1:0] in1,
	input [DATA_WIDTH - 1:0] in2,
	output [DATA_WIDTH - 1:0] out
	);
///////////////////////////////////////////////////////////////
//////////////this code is not complete////////////////////////
///////////////////////////////////////////////////////////////
endmodule
