`timescale 1ns / 1ps


module 
 mem_array_U7_D200 #(parameter
///////////advanced parameters//////////
	DATA_WIDTH 					= 32,
///////////architecture parameters//////
	IFM_SIZE              = 10,                                                
    NUMBER_OF_IFM         = 200,
    NUMBER_OF_UNITS       = 7,
    ADDRESS_SIZE_IFM      = $clog2(IFM_SIZE*IFM_SIZE))

	)(
	input clk,
	input [$clog2($ceil(NUMBER_OF_IFM/NUMBER_OF_UNITS))-1:0] ifm_sel,
	input                        ifm_enable_write_previous,            
	input                        ifm_enable_read_previous, 
	input  [ADDRESS_SIZE_IFM-1:0] ifm_address_write_previous,
	input  [ADDRESS_SIZE_IFM-1:0] ifm_address_read_previous,	

	input [DATA_WIDTH-1:0] data_in_from_previous1,
	input [DATA_WIDTH-1:0] data_in_from_previous2,
	input [DATA_WIDTH-1:0] data_in_from_previous3,
	input [DATA_WIDTH-1:0] data_in_from_previous4,
	input [DATA_WIDTH-1:0] data_in_from_previous5,
	input [DATA_WIDTH-1:0] data_in_from_previous6,
	input [DATA_WIDTH-1:0] data_in_from_previous7,
	output reg [DATA_WIDTH-1:0] data_out_for_previous1,
	output reg [DATA_WIDTH-1:0] data_out_for_previous2,
	output reg [DATA_WIDTH-1:0] data_out_for_previous3,
	output reg [DATA_WIDTH-1:0] data_out_for_previous4,
	output reg [DATA_WIDTH-1:0] data_out_for_previous5,
	output reg [DATA_WIDTH-1:0] data_out_for_previous6,
	output reg [DATA_WIDTH-1:0] data_out_for_previous7,
	input                        ifm_enable_read_A_next,
    input                        ifm_enable_read_B_next,
	input [ADDRESS_SIZE_IFM-1:0] ifm_address_read_A_next,
	input [ADDRESS_SIZE_IFM-1:0] ifm_address_read_B_next,
	output reg [DATA_WIDTH-1:0] data_out_A_for_next1,
	output reg [DATA_WIDTH-1:0] data_out_B_for_next1,
	output reg [DATA_WIDTH-1:0] data_out_A_for_next2,
	output reg [DATA_WIDTH-1:0] data_out_B_for_next2,
	output reg [DATA_WIDTH-1:0] data_out_A_for_next3,
	output reg [DATA_WIDTH-1:0] data_out_B_for_next3,
	output reg [DATA_WIDTH-1:0] data_out_A_for_next4,
	output reg [DATA_WIDTH-1:0] data_out_B_for_next4,
	output reg [DATA_WIDTH-1:0] data_out_A_for_next5,
	output reg [DATA_WIDTH-1:0] data_out_B_for_next5,
	output reg [DATA_WIDTH-1:0] data_out_A_for_next6,
	output reg [DATA_WIDTH-1:0] data_out_B_for_next6,
	output reg [DATA_WIDTH-1:0] data_out_A_for_next7,
	output reg [DATA_WIDTH-1:0] data_out_B_for_next7
	);
	
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem1;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem1;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem2;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem2;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem3;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem3;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem4;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem4;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem5;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem5;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem6;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem6;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem7;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem7;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem8;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem8;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem9;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem9;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem10;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem10;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem11;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem11;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem12;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem12;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem13;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem13;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem14;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem14;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem15;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem15;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem16;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem16;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem17;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem17;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem18;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem18;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem19;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem19;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem20;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem20;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem21;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem21;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem22;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem22;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem23;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem23;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem24;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem24;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem25;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem25;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem26;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem26;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem27;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem27;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem28;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem28;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem29;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem29;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem30;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem30;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem31;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem31;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem32;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem32;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem33;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem33;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem34;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem34;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem35;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem35;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem36;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem36;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem37;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem37;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem38;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem38;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem39;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem39;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem40;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem40;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem41;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem41;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem42;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem42;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem43;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem43;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem44;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem44;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem45;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem45;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem46;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem46;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem47;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem47;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem48;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem48;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem49;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem49;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem50;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem50;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem51;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem51;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem52;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem52;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem53;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem53;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem54;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem54;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem55;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem55;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem56;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem56;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem57;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem57;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem58;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem58;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem59;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem59;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem60;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem60;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem61;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem61;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem62;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem62;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem63;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem63;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem64;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem64;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem65;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem65;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem66;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem66;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem67;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem67;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem68;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem68;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem69;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem69;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem70;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem70;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem71;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem71;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem72;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem72;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem73;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem73;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem74;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem74;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem75;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem75;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem76;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem76;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem77;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem77;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem78;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem78;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem79;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem79;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem80;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem80;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem81;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem81;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem82;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem82;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem83;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem83;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem84;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem84;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem85;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem85;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem86;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem86;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem87;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem87;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem88;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem88;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem89;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem89;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem90;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem90;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem91;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem91;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem92;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem92;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem93;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem93;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem94;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem94;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem95;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem95;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem96;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem96;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem97;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem97;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem98;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem98;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem99;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem99;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem100;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem100;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem101;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem101;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem102;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem102;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem103;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem103;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem104;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem104;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem105;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem105;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem106;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem106;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem107;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem107;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem108;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem108;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem109;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem109;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem110;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem110;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem111;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem111;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem112;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem112;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem113;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem113;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem114;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem114;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem115;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem115;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem116;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem116;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem117;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem117;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem118;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem118;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem119;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem119;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem120;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem120;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem121;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem121;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem122;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem122;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem123;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem123;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem124;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem124;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem125;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem125;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem126;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem126;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem127;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem127;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem128;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem128;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem129;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem129;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem130;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem130;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem131;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem131;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem132;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem132;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem133;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem133;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem134;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem134;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem135;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem135;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem136;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem136;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem137;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem137;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem138;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem138;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem139;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem139;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem140;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem140;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem141;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem141;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem142;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem142;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem143;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem143;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem144;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem144;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem145;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem145;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem146;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem146;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem147;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem147;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem148;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem148;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem149;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem149;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem150;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem150;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem151;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem151;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem152;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem152;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem153;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem153;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem154;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem154;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem155;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem155;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem156;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem156;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem157;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem157;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem158;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem158;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem159;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem159;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem160;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem160;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem161;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem161;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem162;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem162;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem163;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem163;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem164;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem164;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem165;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem165;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem166;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem166;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem167;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem167;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem168;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem168;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem169;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem169;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem170;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem170;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem171;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem171;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem172;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem172;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem173;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem173;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem174;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem174;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem175;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem175;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem176;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem176;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem177;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem177;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem178;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem178;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem179;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem179;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem180;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem180;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem181;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem181;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem182;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem182;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem183;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem183;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem184;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem184;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem185;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem185;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem186;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem186;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem187;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem187;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem188;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem188;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem189;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem189;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem190;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem190;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem191;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem191;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem192;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem192;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem193;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem193;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem194;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem194;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem195;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem195;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem196;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem196;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem197;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem197;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem198;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem198;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem199;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem199;
	wire [DATA_WIDTH-1:0] Data_Output_A_Mem200;
	wire [DATA_WIDTH-1:0] Data_Output_B_Mem200;
	
	wire ifm_enable_write_previous_dMuxOut1;
	wire ifm_enable_read_previous_dMuxOut1;
	wire ifm_enable_read_A_next_dMuxOut1;
	wire ifm_enable_read_B_next_dMuxOut1;
	
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_write_previous_dMuxOut1;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_previous_dMuxOut1;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_A_next_dMuxOut1;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_B_next_dMuxOut1;
	
	
	wire ifm_enable_write_previous_dMuxOut2;
	wire ifm_enable_read_previous_dMuxOut2;
	wire ifm_enable_read_A_next_dMuxOut2;
	wire ifm_enable_read_B_next_dMuxOut2;
	
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_write_previous_dMuxOut2;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_previous_dMuxOut2;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_A_next_dMuxOut2;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_B_next_dMuxOut2;
	
	
	wire ifm_enable_write_previous_dMuxOut3;
	wire ifm_enable_read_previous_dMuxOut3;
	wire ifm_enable_read_A_next_dMuxOut3;
	wire ifm_enable_read_B_next_dMuxOut3;
	
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_write_previous_dMuxOut3;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_previous_dMuxOut3;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_A_next_dMuxOut3;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_B_next_dMuxOut3;
	
	
	wire ifm_enable_write_previous_dMuxOut4;
	wire ifm_enable_read_previous_dMuxOut4;
	wire ifm_enable_read_A_next_dMuxOut4;
	wire ifm_enable_read_B_next_dMuxOut4;
	
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_write_previous_dMuxOut4;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_previous_dMuxOut4;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_A_next_dMuxOut4;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_B_next_dMuxOut4;
	
	
	wire ifm_enable_write_previous_dMuxOut5;
	wire ifm_enable_read_previous_dMuxOut5;
	wire ifm_enable_read_A_next_dMuxOut5;
	wire ifm_enable_read_B_next_dMuxOut5;
	
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_write_previous_dMuxOut5;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_previous_dMuxOut5;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_A_next_dMuxOut5;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_B_next_dMuxOut5;
	
	
	wire ifm_enable_write_previous_dMuxOut6;
	wire ifm_enable_read_previous_dMuxOut6;
	wire ifm_enable_read_A_next_dMuxOut6;
	wire ifm_enable_read_B_next_dMuxOut6;
	
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_write_previous_dMuxOut6;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_previous_dMuxOut6;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_A_next_dMuxOut6;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_B_next_dMuxOut6;
	
	
	wire ifm_enable_write_previous_dMuxOut7;
	wire ifm_enable_read_previous_dMuxOut7;
	wire ifm_enable_read_A_next_dMuxOut7;
	wire ifm_enable_read_B_next_dMuxOut7;
	
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_write_previous_dMuxOut7;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_previous_dMuxOut7;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_A_next_dMuxOut7;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_B_next_dMuxOut7;
	
	
	wire ifm_enable_write_previous_dMuxOut8;
	wire ifm_enable_read_previous_dMuxOut8;
	wire ifm_enable_read_A_next_dMuxOut8;
	wire ifm_enable_read_B_next_dMuxOut8;
	
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_write_previous_dMuxOut8;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_previous_dMuxOut8;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_A_next_dMuxOut8;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_B_next_dMuxOut8;
	
	
	wire ifm_enable_write_previous_dMuxOut9;
	wire ifm_enable_read_previous_dMuxOut9;
	wire ifm_enable_read_A_next_dMuxOut9;
	wire ifm_enable_read_B_next_dMuxOut9;
	
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_write_previous_dMuxOut9;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_previous_dMuxOut9;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_A_next_dMuxOut9;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_B_next_dMuxOut9;
	
	
	wire ifm_enable_write_previous_dMuxOut10;
	wire ifm_enable_read_previous_dMuxOut10;
	wire ifm_enable_read_A_next_dMuxOut10;
	wire ifm_enable_read_B_next_dMuxOut10;
	
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_write_previous_dMuxOut10;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_previous_dMuxOut10;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_A_next_dMuxOut10;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_B_next_dMuxOut10;
	
	
	wire ifm_enable_write_previous_dMuxOut11;
	wire ifm_enable_read_previous_dMuxOut11;
	wire ifm_enable_read_A_next_dMuxOut11;
	wire ifm_enable_read_B_next_dMuxOut11;
	
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_write_previous_dMuxOut11;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_previous_dMuxOut11;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_A_next_dMuxOut11;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_B_next_dMuxOut11;
	
	
	wire ifm_enable_write_previous_dMuxOut12;
	wire ifm_enable_read_previous_dMuxOut12;
	wire ifm_enable_read_A_next_dMuxOut12;
	wire ifm_enable_read_B_next_dMuxOut12;
	
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_write_previous_dMuxOut12;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_previous_dMuxOut12;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_A_next_dMuxOut12;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_B_next_dMuxOut12;
	
	
	wire ifm_enable_write_previous_dMuxOut13;
	wire ifm_enable_read_previous_dMuxOut13;
	wire ifm_enable_read_A_next_dMuxOut13;
	wire ifm_enable_read_B_next_dMuxOut13;
	
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_write_previous_dMuxOut13;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_previous_dMuxOut13;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_A_next_dMuxOut13;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_B_next_dMuxOut13;
	
	
	wire ifm_enable_write_previous_dMuxOut14;
	wire ifm_enable_read_previous_dMuxOut14;
	wire ifm_enable_read_A_next_dMuxOut14;
	wire ifm_enable_read_B_next_dMuxOut14;
	
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_write_previous_dMuxOut14;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_previous_dMuxOut14;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_A_next_dMuxOut14;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_B_next_dMuxOut14;
	
	
	wire ifm_enable_write_previous_dMuxOut15;
	wire ifm_enable_read_previous_dMuxOut15;
	wire ifm_enable_read_A_next_dMuxOut15;
	wire ifm_enable_read_B_next_dMuxOut15;
	
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_write_previous_dMuxOut15;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_previous_dMuxOut15;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_A_next_dMuxOut15;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_B_next_dMuxOut15;
	
	
	wire ifm_enable_write_previous_dMuxOut16;
	wire ifm_enable_read_previous_dMuxOut16;
	wire ifm_enable_read_A_next_dMuxOut16;
	wire ifm_enable_read_B_next_dMuxOut16;
	
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_write_previous_dMuxOut16;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_previous_dMuxOut16;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_A_next_dMuxOut16;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_B_next_dMuxOut16;
	
	
	wire ifm_enable_write_previous_dMuxOut17;
	wire ifm_enable_read_previous_dMuxOut17;
	wire ifm_enable_read_A_next_dMuxOut17;
	wire ifm_enable_read_B_next_dMuxOut17;
	
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_write_previous_dMuxOut17;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_previous_dMuxOut17;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_A_next_dMuxOut17;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_B_next_dMuxOut17;
	
	
	wire ifm_enable_write_previous_dMuxOut18;
	wire ifm_enable_read_previous_dMuxOut18;
	wire ifm_enable_read_A_next_dMuxOut18;
	wire ifm_enable_read_B_next_dMuxOut18;
	
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_write_previous_dMuxOut18;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_previous_dMuxOut18;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_A_next_dMuxOut18;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_B_next_dMuxOut18;
	
	
	wire ifm_enable_write_previous_dMuxOut19;
	wire ifm_enable_read_previous_dMuxOut19;
	wire ifm_enable_read_A_next_dMuxOut19;
	wire ifm_enable_read_B_next_dMuxOut19;
	
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_write_previous_dMuxOut19;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_previous_dMuxOut19;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_A_next_dMuxOut19;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_B_next_dMuxOut19;
	
	
	wire ifm_enable_write_previous_dMuxOut20;
	wire ifm_enable_read_previous_dMuxOut20;
	wire ifm_enable_read_A_next_dMuxOut20;
	wire ifm_enable_read_B_next_dMuxOut20;
	
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_write_previous_dMuxOut20;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_previous_dMuxOut20;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_A_next_dMuxOut20;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_B_next_dMuxOut20;
	
	
	wire ifm_enable_write_previous_dMuxOut21;
	wire ifm_enable_read_previous_dMuxOut21;
	wire ifm_enable_read_A_next_dMuxOut21;
	wire ifm_enable_read_B_next_dMuxOut21;
	
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_write_previous_dMuxOut21;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_previous_dMuxOut21;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_A_next_dMuxOut21;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_B_next_dMuxOut21;
	
	
	wire ifm_enable_write_previous_dMuxOut22;
	wire ifm_enable_read_previous_dMuxOut22;
	wire ifm_enable_read_A_next_dMuxOut22;
	wire ifm_enable_read_B_next_dMuxOut22;
	
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_write_previous_dMuxOut22;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_previous_dMuxOut22;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_A_next_dMuxOut22;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_B_next_dMuxOut22;
	
	
	wire ifm_enable_write_previous_dMuxOut23;
	wire ifm_enable_read_previous_dMuxOut23;
	wire ifm_enable_read_A_next_dMuxOut23;
	wire ifm_enable_read_B_next_dMuxOut23;
	
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_write_previous_dMuxOut23;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_previous_dMuxOut23;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_A_next_dMuxOut23;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_B_next_dMuxOut23;
	
	
	wire ifm_enable_write_previous_dMuxOut24;
	wire ifm_enable_read_previous_dMuxOut24;
	wire ifm_enable_read_A_next_dMuxOut24;
	wire ifm_enable_read_B_next_dMuxOut24;
	
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_write_previous_dMuxOut24;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_previous_dMuxOut24;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_A_next_dMuxOut24;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_B_next_dMuxOut24;
	
	
	wire ifm_enable_write_previous_dMuxOut25;
	wire ifm_enable_read_previous_dMuxOut25;
	wire ifm_enable_read_A_next_dMuxOut25;
	wire ifm_enable_read_B_next_dMuxOut25;
	
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_write_previous_dMuxOut25;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_previous_dMuxOut25;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_A_next_dMuxOut25;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_B_next_dMuxOut25;
	
	
	wire ifm_enable_write_previous_dMuxOut26;
	wire ifm_enable_read_previous_dMuxOut26;
	wire ifm_enable_read_A_next_dMuxOut26;
	wire ifm_enable_read_B_next_dMuxOut26;
	
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_write_previous_dMuxOut26;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_previous_dMuxOut26;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_A_next_dMuxOut26;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_B_next_dMuxOut26;
	
	
	wire ifm_enable_write_previous_dMuxOut27;
	wire ifm_enable_read_previous_dMuxOut27;
	wire ifm_enable_read_A_next_dMuxOut27;
	wire ifm_enable_read_B_next_dMuxOut27;
	
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_write_previous_dMuxOut27;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_previous_dMuxOut27;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_A_next_dMuxOut27;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_B_next_dMuxOut27;
	
	
	wire ifm_enable_write_previous_dMuxOut28;
	wire ifm_enable_read_previous_dMuxOut28;
	wire ifm_enable_read_A_next_dMuxOut28;
	wire ifm_enable_read_B_next_dMuxOut28;
	
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_write_previous_dMuxOut28;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_previous_dMuxOut28;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_A_next_dMuxOut28;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_B_next_dMuxOut28;
	
	
	wire ifm_enable_write_previous_dMuxOut29;
	wire ifm_enable_read_previous_dMuxOut29;
	wire ifm_enable_read_A_next_dMuxOut29;
	wire ifm_enable_read_B_next_dMuxOut29;
	
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_write_previous_dMuxOut29;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_previous_dMuxOut29;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_A_next_dMuxOut29;
	wire [ADDRESS_SIZE_IFM-1:0] ifm_address_read_B_next_dMuxOut29;
	
	demux_1_to_29 d0(
	.din(ifm_enable_write_previous),
	.sel(ifm_sel),
	.dout_1(ifm_enable_write_previous_dMuxOut1),
	.dout_2(ifm_enable_write_previous_dMuxOut2),
	.dout_3(ifm_enable_write_previous_dMuxOut3),
	.dout_4(ifm_enable_write_previous_dMuxOut4),
	.dout_5(ifm_enable_write_previous_dMuxOut5),
	.dout_6(ifm_enable_write_previous_dMuxOut6),
	.dout_7(ifm_enable_write_previous_dMuxOut7),
	.dout_8(ifm_enable_write_previous_dMuxOut8),
	.dout_9(ifm_enable_write_previous_dMuxOut9),
	.dout_10(ifm_enable_write_previous_dMuxOut10),
	.dout_11(ifm_enable_write_previous_dMuxOut11),
	.dout_12(ifm_enable_write_previous_dMuxOut12),
	.dout_13(ifm_enable_write_previous_dMuxOut13),
	.dout_14(ifm_enable_write_previous_dMuxOut14),
	.dout_15(ifm_enable_write_previous_dMuxOut15),
	.dout_16(ifm_enable_write_previous_dMuxOut16),
	.dout_17(ifm_enable_write_previous_dMuxOut17),
	.dout_18(ifm_enable_write_previous_dMuxOut18),
	.dout_19(ifm_enable_write_previous_dMuxOut19),
	.dout_20(ifm_enable_write_previous_dMuxOut20),
	.dout_21(ifm_enable_write_previous_dMuxOut21),
	.dout_22(ifm_enable_write_previous_dMuxOut22),
	.dout_23(ifm_enable_write_previous_dMuxOut23),
	.dout_24(ifm_enable_write_previous_dMuxOut24),
	.dout_25(ifm_enable_write_previous_dMuxOut25),
	.dout_26(ifm_enable_write_previous_dMuxOut26),
	.dout_27(ifm_enable_write_previous_dMuxOut27),
	.dout_28(ifm_enable_write_previous_dMuxOut28),
	.dout_29(ifm_enable_write_previous_dMuxOut29)
	);

	demux_1_to_29 d1(
	.din(ifm_enable_read_previous),
	.sel(ifm_sel),
	.dout_1(ifm_enable_read_previous_dMuxOut1),
	.dout_2(ifm_enable_read_previous_dMuxOut2),
	.dout_3(ifm_enable_read_previous_dMuxOut3),
	.dout_4(ifm_enable_read_previous_dMuxOut4),
	.dout_5(ifm_enable_read_previous_dMuxOut5),
	.dout_6(ifm_enable_read_previous_dMuxOut6),
	.dout_7(ifm_enable_read_previous_dMuxOut7),
	.dout_8(ifm_enable_read_previous_dMuxOut8),
	.dout_9(ifm_enable_read_previous_dMuxOut9),
	.dout_10(ifm_enable_read_previous_dMuxOut10),
	.dout_11(ifm_enable_read_previous_dMuxOut11),
	.dout_12(ifm_enable_read_previous_dMuxOut12),
	.dout_13(ifm_enable_read_previous_dMuxOut13),
	.dout_14(ifm_enable_read_previous_dMuxOut14),
	.dout_15(ifm_enable_read_previous_dMuxOut15),
	.dout_16(ifm_enable_read_previous_dMuxOut16),
	.dout_17(ifm_enable_read_previous_dMuxOut17),
	.dout_18(ifm_enable_read_previous_dMuxOut18),
	.dout_19(ifm_enable_read_previous_dMuxOut19),
	.dout_20(ifm_enable_read_previous_dMuxOut20),
	.dout_21(ifm_enable_read_previous_dMuxOut21),
	.dout_22(ifm_enable_read_previous_dMuxOut22),
	.dout_23(ifm_enable_read_previous_dMuxOut23),
	.dout_24(ifm_enable_read_previous_dMuxOut24),
	.dout_25(ifm_enable_read_previous_dMuxOut25),
	.dout_26(ifm_enable_read_previous_dMuxOut26),
	.dout_27(ifm_enable_read_previous_dMuxOut27),
	.dout_28(ifm_enable_read_previous_dMuxOut28),
	.dout_29(ifm_enable_read_previous_dMuxOut29)
	);

	demux_1_to_29 d2(
	.din(ifm_enable_read_B_next),
	.sel(ifm_sel),
	.dout_1(ifm_enable_read_B_next_dMuxOut1),
	.dout_2(ifm_enable_read_B_next_dMuxOut2),
	.dout_3(ifm_enable_read_B_next_dMuxOut3),
	.dout_4(ifm_enable_read_B_next_dMuxOut4),
	.dout_5(ifm_enable_read_B_next_dMuxOut5),
	.dout_6(ifm_enable_read_B_next_dMuxOut6),
	.dout_7(ifm_enable_read_B_next_dMuxOut7),
	.dout_8(ifm_enable_read_B_next_dMuxOut8),
	.dout_9(ifm_enable_read_B_next_dMuxOut9),
	.dout_10(ifm_enable_read_B_next_dMuxOut10),
	.dout_11(ifm_enable_read_B_next_dMuxOut11),
	.dout_12(ifm_enable_read_B_next_dMuxOut12),
	.dout_13(ifm_enable_read_B_next_dMuxOut13),
	.dout_14(ifm_enable_read_B_next_dMuxOut14),
	.dout_15(ifm_enable_read_B_next_dMuxOut15),
	.dout_16(ifm_enable_read_B_next_dMuxOut16),
	.dout_17(ifm_enable_read_B_next_dMuxOut17),
	.dout_18(ifm_enable_read_B_next_dMuxOut18),
	.dout_19(ifm_enable_read_B_next_dMuxOut19),
	.dout_20(ifm_enable_read_B_next_dMuxOut20),
	.dout_21(ifm_enable_read_B_next_dMuxOut21),
	.dout_22(ifm_enable_read_B_next_dMuxOut22),
	.dout_23(ifm_enable_read_B_next_dMuxOut23),
	.dout_24(ifm_enable_read_B_next_dMuxOut24),
	.dout_25(ifm_enable_read_B_next_dMuxOut25),
	.dout_26(ifm_enable_read_B_next_dMuxOut26),
	.dout_27(ifm_enable_read_B_next_dMuxOut27),
	.dout_28(ifm_enable_read_B_next_dMuxOut28),
	.dout_29(ifm_enable_read_B_next_dMuxOut29)
	);

	demux_1_to_29 d3(
	.din(ifm_enable_write_previous),
	.sel(ifm_sel),
	.dout_1(ifm_enable_write_previous_dMuxOut1),
	.dout_2(ifm_enable_write_previous_dMuxOut2),
	.dout_3(ifm_enable_write_previous_dMuxOut3),
	.dout_4(ifm_enable_write_previous_dMuxOut4),
	.dout_5(ifm_enable_write_previous_dMuxOut5),
	.dout_6(ifm_enable_write_previous_dMuxOut6),
	.dout_7(ifm_enable_write_previous_dMuxOut7),
	.dout_8(ifm_enable_write_previous_dMuxOut8),
	.dout_9(ifm_enable_write_previous_dMuxOut9),
	.dout_10(ifm_enable_write_previous_dMuxOut10),
	.dout_11(ifm_enable_write_previous_dMuxOut11),
	.dout_12(ifm_enable_write_previous_dMuxOut12),
	.dout_13(ifm_enable_write_previous_dMuxOut13),
	.dout_14(ifm_enable_write_previous_dMuxOut14),
	.dout_15(ifm_enable_write_previous_dMuxOut15),
	.dout_16(ifm_enable_write_previous_dMuxOut16),
	.dout_17(ifm_enable_write_previous_dMuxOut17),
	.dout_18(ifm_enable_write_previous_dMuxOut18),
	.dout_19(ifm_enable_write_previous_dMuxOut19),
	.dout_20(ifm_enable_write_previous_dMuxOut20),
	.dout_21(ifm_enable_write_previous_dMuxOut21),
	.dout_22(ifm_enable_write_previous_dMuxOut22),
	.dout_23(ifm_enable_write_previous_dMuxOut23),
	.dout_24(ifm_enable_write_previous_dMuxOut24),
	.dout_25(ifm_enable_write_previous_dMuxOut25),
	.dout_26(ifm_enable_write_previous_dMuxOut26),
	.dout_27(ifm_enable_write_previous_dMuxOut27),
	.dout_28(ifm_enable_write_previous_dMuxOut28),
	.dout_29(ifm_enable_write_previous_dMuxOut29)
	);

	demux_1_to_29_7bits d4(
	.din(ifm_address_write_previous),
	.sel(ifm_sel),
	.dout_1(ifm_address_write_previous_dMuxOut1),
	.dout_2(ifm_address_write_previous_dMuxOut2),
	.dout_3(ifm_address_write_previous_dMuxOut3),
	.dout_4(ifm_address_write_previous_dMuxOut4),
	.dout_5(ifm_address_write_previous_dMuxOut5),
	.dout_6(ifm_address_write_previous_dMuxOut6),
	.dout_7(ifm_address_write_previous_dMuxOut7),
	.dout_8(ifm_address_write_previous_dMuxOut8),
	.dout_9(ifm_address_write_previous_dMuxOut9),
	.dout_10(ifm_address_write_previous_dMuxOut10),
	.dout_11(ifm_address_write_previous_dMuxOut11),
	.dout_12(ifm_address_write_previous_dMuxOut12),
	.dout_13(ifm_address_write_previous_dMuxOut13),
	.dout_14(ifm_address_write_previous_dMuxOut14),
	.dout_15(ifm_address_write_previous_dMuxOut15),
	.dout_16(ifm_address_write_previous_dMuxOut16),
	.dout_17(ifm_address_write_previous_dMuxOut17),
	.dout_18(ifm_address_write_previous_dMuxOut18),
	.dout_19(ifm_address_write_previous_dMuxOut19),
	.dout_20(ifm_address_write_previous_dMuxOut20),
	.dout_21(ifm_address_write_previous_dMuxOut21),
	.dout_22(ifm_address_write_previous_dMuxOut22),
	.dout_23(ifm_address_write_previous_dMuxOut23),
	.dout_24(ifm_address_write_previous_dMuxOut24),
	.dout_25(ifm_address_write_previous_dMuxOut25),
	.dout_26(ifm_address_write_previous_dMuxOut26),
	.dout_27(ifm_address_write_previous_dMuxOut27),
	.dout_28(ifm_address_write_previous_dMuxOut28),
	.dout_29(ifm_address_write_previous_dMuxOut29)
	);

	demux_1_to_29_7bits d5(
	.din(ifm_address_read_previous),
	.sel(ifm_sel),
	.dout_1(ifm_address_read_previous_dMuxOut1),
	.dout_2(ifm_address_read_previous_dMuxOut2),
	.dout_3(ifm_address_read_previous_dMuxOut3),
	.dout_4(ifm_address_read_previous_dMuxOut4),
	.dout_5(ifm_address_read_previous_dMuxOut5),
	.dout_6(ifm_address_read_previous_dMuxOut6),
	.dout_7(ifm_address_read_previous_dMuxOut7),
	.dout_8(ifm_address_read_previous_dMuxOut8),
	.dout_9(ifm_address_read_previous_dMuxOut9),
	.dout_10(ifm_address_read_previous_dMuxOut10),
	.dout_11(ifm_address_read_previous_dMuxOut11),
	.dout_12(ifm_address_read_previous_dMuxOut12),
	.dout_13(ifm_address_read_previous_dMuxOut13),
	.dout_14(ifm_address_read_previous_dMuxOut14),
	.dout_15(ifm_address_read_previous_dMuxOut15),
	.dout_16(ifm_address_read_previous_dMuxOut16),
	.dout_17(ifm_address_read_previous_dMuxOut17),
	.dout_18(ifm_address_read_previous_dMuxOut18),
	.dout_19(ifm_address_read_previous_dMuxOut19),
	.dout_20(ifm_address_read_previous_dMuxOut20),
	.dout_21(ifm_address_read_previous_dMuxOut21),
	.dout_22(ifm_address_read_previous_dMuxOut22),
	.dout_23(ifm_address_read_previous_dMuxOut23),
	.dout_24(ifm_address_read_previous_dMuxOut24),
	.dout_25(ifm_address_read_previous_dMuxOut25),
	.dout_26(ifm_address_read_previous_dMuxOut26),
	.dout_27(ifm_address_read_previous_dMuxOut27),
	.dout_28(ifm_address_read_previous_dMuxOut28),
	.dout_29(ifm_address_read_previous_dMuxOut29)
	);

	demux_1_to_29_7bits d6(
	.din(ifm_address_read_A_next),
	.sel(ifm_sel),
	.dout_1(ifm_address_read_A_next_dMuxOut1),
	.dout_2(ifm_address_read_A_next_dMuxOut2),
	.dout_3(ifm_address_read_A_next_dMuxOut3),
	.dout_4(ifm_address_read_A_next_dMuxOut4),
	.dout_5(ifm_address_read_A_next_dMuxOut5),
	.dout_6(ifm_address_read_A_next_dMuxOut6),
	.dout_7(ifm_address_read_A_next_dMuxOut7),
	.dout_8(ifm_address_read_A_next_dMuxOut8),
	.dout_9(ifm_address_read_A_next_dMuxOut9),
	.dout_10(ifm_address_read_A_next_dMuxOut10),
	.dout_11(ifm_address_read_A_next_dMuxOut11),
	.dout_12(ifm_address_read_A_next_dMuxOut12),
	.dout_13(ifm_address_read_A_next_dMuxOut13),
	.dout_14(ifm_address_read_A_next_dMuxOut14),
	.dout_15(ifm_address_read_A_next_dMuxOut15),
	.dout_16(ifm_address_read_A_next_dMuxOut16),
	.dout_17(ifm_address_read_A_next_dMuxOut17),
	.dout_18(ifm_address_read_A_next_dMuxOut18),
	.dout_19(ifm_address_read_A_next_dMuxOut19),
	.dout_20(ifm_address_read_A_next_dMuxOut20),
	.dout_21(ifm_address_read_A_next_dMuxOut21),
	.dout_22(ifm_address_read_A_next_dMuxOut22),
	.dout_23(ifm_address_read_A_next_dMuxOut23),
	.dout_24(ifm_address_read_A_next_dMuxOut24),
	.dout_25(ifm_address_read_A_next_dMuxOut25),
	.dout_26(ifm_address_read_A_next_dMuxOut26),
	.dout_27(ifm_address_read_A_next_dMuxOut27),
	.dout_28(ifm_address_read_A_next_dMuxOut28),
	.dout_29(ifm_address_read_A_next_dMuxOut29)
	);

	demux_1_to_29_7bits d7(
	.din(ifm_address_read_B_next),
	.sel(ifm_sel),
	.dout_1(ifm_address_read_B_next_dMuxOut1),
	.dout_2(ifm_address_read_B_next_dMuxOut2),
	.dout_3(ifm_address_read_B_next_dMuxOut3),
	.dout_4(ifm_address_read_B_next_dMuxOut4),
	.dout_5(ifm_address_read_B_next_dMuxOut5),
	.dout_6(ifm_address_read_B_next_dMuxOut6),
	.dout_7(ifm_address_read_B_next_dMuxOut7),
	.dout_8(ifm_address_read_B_next_dMuxOut8),
	.dout_9(ifm_address_read_B_next_dMuxOut9),
	.dout_10(ifm_address_read_B_next_dMuxOut10),
	.dout_11(ifm_address_read_B_next_dMuxOut11),
	.dout_12(ifm_address_read_B_next_dMuxOut12),
	.dout_13(ifm_address_read_B_next_dMuxOut13),
	.dout_14(ifm_address_read_B_next_dMuxOut14),
	.dout_15(ifm_address_read_B_next_dMuxOut15),
	.dout_16(ifm_address_read_B_next_dMuxOut16),
	.dout_17(ifm_address_read_B_next_dMuxOut17),
	.dout_18(ifm_address_read_B_next_dMuxOut18),
	.dout_19(ifm_address_read_B_next_dMuxOut19),
	.dout_20(ifm_address_read_B_next_dMuxOut20),
	.dout_21(ifm_address_read_B_next_dMuxOut21),
	.dout_22(ifm_address_read_B_next_dMuxOut22),
	.dout_23(ifm_address_read_B_next_dMuxOut23),
	.dout_24(ifm_address_read_B_next_dMuxOut24),
	.dout_25(ifm_address_read_B_next_dMuxOut25),
	.dout_26(ifm_address_read_B_next_dMuxOut26),
	.dout_27(ifm_address_read_B_next_dMuxOut27),
	.dout_28(ifm_address_read_B_next_dMuxOut28),
	.dout_29(ifm_address_read_B_next_dMuxOut29)
	);

	
    always @*
    begin

        case(ifm_sel)
		5'd0:
		begin
			data_out_for_previous1 = Data_Output_B_Mem1;
			data_out_for_previous2 = Data_Output_B_Mem2;
			data_out_for_previous3 = Data_Output_B_Mem3;
			data_out_for_previous4 = Data_Output_B_Mem4;
			data_out_for_previous5 = Data_Output_B_Mem5;
			data_out_for_previous6 = Data_Output_B_Mem6;
			data_out_for_previous7 = Data_Output_B_Mem7;
		
			data_out_A_for_next1 = Data_Output_A_Mem197;
			data_out_B_for_next1 = Data_Output_B_Mem197;
		
			data_out_A_for_next2 = Data_Output_A_Mem198;
			data_out_B_for_next2 = Data_Output_B_Mem198;
		
			data_out_A_for_next3 = Data_Output_A_Mem199;
			data_out_B_for_next3 = Data_Output_B_Mem199;
		
			data_out_A_for_next4 = Data_Output_A_Mem200;
			data_out_B_for_next4 = Data_Output_B_Mem200;
		
			data_out_A_for_next5 = 0;
			data_out_B_for_next5 = 0;
		
			data_out_A_for_next6 = 0;
			data_out_B_for_next6 = 0;
		
			data_out_A_for_next7 = 0;
			data_out_B_for_next7 = 0;
		end
		5'd1:
		begin
			data_out_for_previous1 = Data_Output_B_Mem8;
			data_out_for_previous2 = Data_Output_B_Mem9;
			data_out_for_previous3 = Data_Output_B_Mem10;
			data_out_for_previous4 = Data_Output_B_Mem11;
			data_out_for_previous5 = Data_Output_B_Mem12;
			data_out_for_previous6 = Data_Output_B_Mem13;
			data_out_for_previous7 = Data_Output_B_Mem14;
		
			data_out_A_for_next1 = Data_Output_A_Mem1;
			data_out_B_for_next1 = Data_Output_B_Mem1;
		
			data_out_A_for_next2 = Data_Output_A_Mem2;
			data_out_B_for_next2 = Data_Output_B_Mem2;
		
			data_out_A_for_next3 = Data_Output_A_Mem3;
			data_out_B_for_next3 = Data_Output_B_Mem3;
		
			data_out_A_for_next4 = Data_Output_A_Mem4;
			data_out_B_for_next4 = Data_Output_B_Mem4;
		
			data_out_A_for_next5 = Data_Output_A_Mem5;
			data_out_B_for_next5 = Data_Output_B_Mem5;
		
			data_out_A_for_next6 = Data_Output_A_Mem6;
			data_out_B_for_next6 = Data_Output_B_Mem6;
		
			data_out_A_for_next7 = Data_Output_A_Mem7;
			data_out_B_for_next7 = Data_Output_B_Mem7;
		end
		5'd2:
		begin
			data_out_for_previous1 = Data_Output_B_Mem15;
			data_out_for_previous2 = Data_Output_B_Mem16;
			data_out_for_previous3 = Data_Output_B_Mem17;
			data_out_for_previous4 = Data_Output_B_Mem18;
			data_out_for_previous5 = Data_Output_B_Mem19;
			data_out_for_previous6 = Data_Output_B_Mem20;
			data_out_for_previous7 = Data_Output_B_Mem21;
		
			data_out_A_for_next1 = Data_Output_A_Mem8;
			data_out_B_for_next1 = Data_Output_B_Mem8;
		
			data_out_A_for_next2 = Data_Output_A_Mem9;
			data_out_B_for_next2 = Data_Output_B_Mem9;
		
			data_out_A_for_next3 = Data_Output_A_Mem10;
			data_out_B_for_next3 = Data_Output_B_Mem10;
		
			data_out_A_for_next4 = Data_Output_A_Mem11;
			data_out_B_for_next4 = Data_Output_B_Mem11;
		
			data_out_A_for_next5 = Data_Output_A_Mem12;
			data_out_B_for_next5 = Data_Output_B_Mem12;
		
			data_out_A_for_next6 = Data_Output_A_Mem13;
			data_out_B_for_next6 = Data_Output_B_Mem13;
		
			data_out_A_for_next7 = Data_Output_A_Mem14;
			data_out_B_for_next7 = Data_Output_B_Mem14;
		end
		5'd3:
		begin
			data_out_for_previous1 = Data_Output_B_Mem22;
			data_out_for_previous2 = Data_Output_B_Mem23;
			data_out_for_previous3 = Data_Output_B_Mem24;
			data_out_for_previous4 = Data_Output_B_Mem25;
			data_out_for_previous5 = Data_Output_B_Mem26;
			data_out_for_previous6 = Data_Output_B_Mem27;
			data_out_for_previous7 = Data_Output_B_Mem28;
		
			data_out_A_for_next1 = Data_Output_A_Mem15;
			data_out_B_for_next1 = Data_Output_B_Mem15;
		
			data_out_A_for_next2 = Data_Output_A_Mem16;
			data_out_B_for_next2 = Data_Output_B_Mem16;
		
			data_out_A_for_next3 = Data_Output_A_Mem17;
			data_out_B_for_next3 = Data_Output_B_Mem17;
		
			data_out_A_for_next4 = Data_Output_A_Mem18;
			data_out_B_for_next4 = Data_Output_B_Mem18;
		
			data_out_A_for_next5 = Data_Output_A_Mem19;
			data_out_B_for_next5 = Data_Output_B_Mem19;
		
			data_out_A_for_next6 = Data_Output_A_Mem20;
			data_out_B_for_next6 = Data_Output_B_Mem20;
		
			data_out_A_for_next7 = Data_Output_A_Mem21;
			data_out_B_for_next7 = Data_Output_B_Mem21;
		end
		5'd4:
		begin
			data_out_for_previous1 = Data_Output_B_Mem29;
			data_out_for_previous2 = Data_Output_B_Mem30;
			data_out_for_previous3 = Data_Output_B_Mem31;
			data_out_for_previous4 = Data_Output_B_Mem32;
			data_out_for_previous5 = Data_Output_B_Mem33;
			data_out_for_previous6 = Data_Output_B_Mem34;
			data_out_for_previous7 = Data_Output_B_Mem35;
		
			data_out_A_for_next1 = Data_Output_A_Mem22;
			data_out_B_for_next1 = Data_Output_B_Mem22;
		
			data_out_A_for_next2 = Data_Output_A_Mem23;
			data_out_B_for_next2 = Data_Output_B_Mem23;
		
			data_out_A_for_next3 = Data_Output_A_Mem24;
			data_out_B_for_next3 = Data_Output_B_Mem24;
		
			data_out_A_for_next4 = Data_Output_A_Mem25;
			data_out_B_for_next4 = Data_Output_B_Mem25;
		
			data_out_A_for_next5 = Data_Output_A_Mem26;
			data_out_B_for_next5 = Data_Output_B_Mem26;
		
			data_out_A_for_next6 = Data_Output_A_Mem27;
			data_out_B_for_next6 = Data_Output_B_Mem27;
		
			data_out_A_for_next7 = Data_Output_A_Mem28;
			data_out_B_for_next7 = Data_Output_B_Mem28;
		end
		5'd5:
		begin
			data_out_for_previous1 = Data_Output_B_Mem36;
			data_out_for_previous2 = Data_Output_B_Mem37;
			data_out_for_previous3 = Data_Output_B_Mem38;
			data_out_for_previous4 = Data_Output_B_Mem39;
			data_out_for_previous5 = Data_Output_B_Mem40;
			data_out_for_previous6 = Data_Output_B_Mem41;
			data_out_for_previous7 = Data_Output_B_Mem42;
		
			data_out_A_for_next1 = Data_Output_A_Mem29;
			data_out_B_for_next1 = Data_Output_B_Mem29;
		
			data_out_A_for_next2 = Data_Output_A_Mem30;
			data_out_B_for_next2 = Data_Output_B_Mem30;
		
			data_out_A_for_next3 = Data_Output_A_Mem31;
			data_out_B_for_next3 = Data_Output_B_Mem31;
		
			data_out_A_for_next4 = Data_Output_A_Mem32;
			data_out_B_for_next4 = Data_Output_B_Mem32;
		
			data_out_A_for_next5 = Data_Output_A_Mem33;
			data_out_B_for_next5 = Data_Output_B_Mem33;
		
			data_out_A_for_next6 = Data_Output_A_Mem34;
			data_out_B_for_next6 = Data_Output_B_Mem34;
		
			data_out_A_for_next7 = Data_Output_A_Mem35;
			data_out_B_for_next7 = Data_Output_B_Mem35;
		end
		5'd6:
		begin
			data_out_for_previous1 = Data_Output_B_Mem43;
			data_out_for_previous2 = Data_Output_B_Mem44;
			data_out_for_previous3 = Data_Output_B_Mem45;
			data_out_for_previous4 = Data_Output_B_Mem46;
			data_out_for_previous5 = Data_Output_B_Mem47;
			data_out_for_previous6 = Data_Output_B_Mem48;
			data_out_for_previous7 = Data_Output_B_Mem49;
		
			data_out_A_for_next1 = Data_Output_A_Mem36;
			data_out_B_for_next1 = Data_Output_B_Mem36;
		
			data_out_A_for_next2 = Data_Output_A_Mem37;
			data_out_B_for_next2 = Data_Output_B_Mem37;
		
			data_out_A_for_next3 = Data_Output_A_Mem38;
			data_out_B_for_next3 = Data_Output_B_Mem38;
		
			data_out_A_for_next4 = Data_Output_A_Mem39;
			data_out_B_for_next4 = Data_Output_B_Mem39;
		
			data_out_A_for_next5 = Data_Output_A_Mem40;
			data_out_B_for_next5 = Data_Output_B_Mem40;
		
			data_out_A_for_next6 = Data_Output_A_Mem41;
			data_out_B_for_next6 = Data_Output_B_Mem41;
		
			data_out_A_for_next7 = Data_Output_A_Mem42;
			data_out_B_for_next7 = Data_Output_B_Mem42;
		end
		5'd7:
		begin
			data_out_for_previous1 = Data_Output_B_Mem50;
			data_out_for_previous2 = Data_Output_B_Mem51;
			data_out_for_previous3 = Data_Output_B_Mem52;
			data_out_for_previous4 = Data_Output_B_Mem53;
			data_out_for_previous5 = Data_Output_B_Mem54;
			data_out_for_previous6 = Data_Output_B_Mem55;
			data_out_for_previous7 = Data_Output_B_Mem56;
		
			data_out_A_for_next1 = Data_Output_A_Mem43;
			data_out_B_for_next1 = Data_Output_B_Mem43;
		
			data_out_A_for_next2 = Data_Output_A_Mem44;
			data_out_B_for_next2 = Data_Output_B_Mem44;
		
			data_out_A_for_next3 = Data_Output_A_Mem45;
			data_out_B_for_next3 = Data_Output_B_Mem45;
		
			data_out_A_for_next4 = Data_Output_A_Mem46;
			data_out_B_for_next4 = Data_Output_B_Mem46;
		
			data_out_A_for_next5 = Data_Output_A_Mem47;
			data_out_B_for_next5 = Data_Output_B_Mem47;
		
			data_out_A_for_next6 = Data_Output_A_Mem48;
			data_out_B_for_next6 = Data_Output_B_Mem48;
		
			data_out_A_for_next7 = Data_Output_A_Mem49;
			data_out_B_for_next7 = Data_Output_B_Mem49;
		end
		5'd8:
		begin
			data_out_for_previous1 = Data_Output_B_Mem57;
			data_out_for_previous2 = Data_Output_B_Mem58;
			data_out_for_previous3 = Data_Output_B_Mem59;
			data_out_for_previous4 = Data_Output_B_Mem60;
			data_out_for_previous5 = Data_Output_B_Mem61;
			data_out_for_previous6 = Data_Output_B_Mem62;
			data_out_for_previous7 = Data_Output_B_Mem63;
		
			data_out_A_for_next1 = Data_Output_A_Mem50;
			data_out_B_for_next1 = Data_Output_B_Mem50;
		
			data_out_A_for_next2 = Data_Output_A_Mem51;
			data_out_B_for_next2 = Data_Output_B_Mem51;
		
			data_out_A_for_next3 = Data_Output_A_Mem52;
			data_out_B_for_next3 = Data_Output_B_Mem52;
		
			data_out_A_for_next4 = Data_Output_A_Mem53;
			data_out_B_for_next4 = Data_Output_B_Mem53;
		
			data_out_A_for_next5 = Data_Output_A_Mem54;
			data_out_B_for_next5 = Data_Output_B_Mem54;
		
			data_out_A_for_next6 = Data_Output_A_Mem55;
			data_out_B_for_next6 = Data_Output_B_Mem55;
		
			data_out_A_for_next7 = Data_Output_A_Mem56;
			data_out_B_for_next7 = Data_Output_B_Mem56;
		end
		5'd9:
		begin
			data_out_for_previous1 = Data_Output_B_Mem64;
			data_out_for_previous2 = Data_Output_B_Mem65;
			data_out_for_previous3 = Data_Output_B_Mem66;
			data_out_for_previous4 = Data_Output_B_Mem67;
			data_out_for_previous5 = Data_Output_B_Mem68;
			data_out_for_previous6 = Data_Output_B_Mem69;
			data_out_for_previous7 = Data_Output_B_Mem70;
		
			data_out_A_for_next1 = Data_Output_A_Mem57;
			data_out_B_for_next1 = Data_Output_B_Mem57;
		
			data_out_A_for_next2 = Data_Output_A_Mem58;
			data_out_B_for_next2 = Data_Output_B_Mem58;
		
			data_out_A_for_next3 = Data_Output_A_Mem59;
			data_out_B_for_next3 = Data_Output_B_Mem59;
		
			data_out_A_for_next4 = Data_Output_A_Mem60;
			data_out_B_for_next4 = Data_Output_B_Mem60;
		
			data_out_A_for_next5 = Data_Output_A_Mem61;
			data_out_B_for_next5 = Data_Output_B_Mem61;
		
			data_out_A_for_next6 = Data_Output_A_Mem62;
			data_out_B_for_next6 = Data_Output_B_Mem62;
		
			data_out_A_for_next7 = Data_Output_A_Mem63;
			data_out_B_for_next7 = Data_Output_B_Mem63;
		end
		5'd10:
		begin
			data_out_for_previous1 = Data_Output_B_Mem71;
			data_out_for_previous2 = Data_Output_B_Mem72;
			data_out_for_previous3 = Data_Output_B_Mem73;
			data_out_for_previous4 = Data_Output_B_Mem74;
			data_out_for_previous5 = Data_Output_B_Mem75;
			data_out_for_previous6 = Data_Output_B_Mem76;
			data_out_for_previous7 = Data_Output_B_Mem77;
		
			data_out_A_for_next1 = Data_Output_A_Mem64;
			data_out_B_for_next1 = Data_Output_B_Mem64;
		
			data_out_A_for_next2 = Data_Output_A_Mem65;
			data_out_B_for_next2 = Data_Output_B_Mem65;
		
			data_out_A_for_next3 = Data_Output_A_Mem66;
			data_out_B_for_next3 = Data_Output_B_Mem66;
		
			data_out_A_for_next4 = Data_Output_A_Mem67;
			data_out_B_for_next4 = Data_Output_B_Mem67;
		
			data_out_A_for_next5 = Data_Output_A_Mem68;
			data_out_B_for_next5 = Data_Output_B_Mem68;
		
			data_out_A_for_next6 = Data_Output_A_Mem69;
			data_out_B_for_next6 = Data_Output_B_Mem69;
		
			data_out_A_for_next7 = Data_Output_A_Mem70;
			data_out_B_for_next7 = Data_Output_B_Mem70;
		end
		5'd11:
		begin
			data_out_for_previous1 = Data_Output_B_Mem78;
			data_out_for_previous2 = Data_Output_B_Mem79;
			data_out_for_previous3 = Data_Output_B_Mem80;
			data_out_for_previous4 = Data_Output_B_Mem81;
			data_out_for_previous5 = Data_Output_B_Mem82;
			data_out_for_previous6 = Data_Output_B_Mem83;
			data_out_for_previous7 = Data_Output_B_Mem84;
		
			data_out_A_for_next1 = Data_Output_A_Mem71;
			data_out_B_for_next1 = Data_Output_B_Mem71;
		
			data_out_A_for_next2 = Data_Output_A_Mem72;
			data_out_B_for_next2 = Data_Output_B_Mem72;
		
			data_out_A_for_next3 = Data_Output_A_Mem73;
			data_out_B_for_next3 = Data_Output_B_Mem73;
		
			data_out_A_for_next4 = Data_Output_A_Mem74;
			data_out_B_for_next4 = Data_Output_B_Mem74;
		
			data_out_A_for_next5 = Data_Output_A_Mem75;
			data_out_B_for_next5 = Data_Output_B_Mem75;
		
			data_out_A_for_next6 = Data_Output_A_Mem76;
			data_out_B_for_next6 = Data_Output_B_Mem76;
		
			data_out_A_for_next7 = Data_Output_A_Mem77;
			data_out_B_for_next7 = Data_Output_B_Mem77;
		end
		5'd12:
		begin
			data_out_for_previous1 = Data_Output_B_Mem85;
			data_out_for_previous2 = Data_Output_B_Mem86;
			data_out_for_previous3 = Data_Output_B_Mem87;
			data_out_for_previous4 = Data_Output_B_Mem88;
			data_out_for_previous5 = Data_Output_B_Mem89;
			data_out_for_previous6 = Data_Output_B_Mem90;
			data_out_for_previous7 = Data_Output_B_Mem91;
		
			data_out_A_for_next1 = Data_Output_A_Mem78;
			data_out_B_for_next1 = Data_Output_B_Mem78;
		
			data_out_A_for_next2 = Data_Output_A_Mem79;
			data_out_B_for_next2 = Data_Output_B_Mem79;
		
			data_out_A_for_next3 = Data_Output_A_Mem80;
			data_out_B_for_next3 = Data_Output_B_Mem80;
		
			data_out_A_for_next4 = Data_Output_A_Mem81;
			data_out_B_for_next4 = Data_Output_B_Mem81;
		
			data_out_A_for_next5 = Data_Output_A_Mem82;
			data_out_B_for_next5 = Data_Output_B_Mem82;
		
			data_out_A_for_next6 = Data_Output_A_Mem83;
			data_out_B_for_next6 = Data_Output_B_Mem83;
		
			data_out_A_for_next7 = Data_Output_A_Mem84;
			data_out_B_for_next7 = Data_Output_B_Mem84;
		end
		5'd13:
		begin
			data_out_for_previous1 = Data_Output_B_Mem92;
			data_out_for_previous2 = Data_Output_B_Mem93;
			data_out_for_previous3 = Data_Output_B_Mem94;
			data_out_for_previous4 = Data_Output_B_Mem95;
			data_out_for_previous5 = Data_Output_B_Mem96;
			data_out_for_previous6 = Data_Output_B_Mem97;
			data_out_for_previous7 = Data_Output_B_Mem98;
		
			data_out_A_for_next1 = Data_Output_A_Mem85;
			data_out_B_for_next1 = Data_Output_B_Mem85;
		
			data_out_A_for_next2 = Data_Output_A_Mem86;
			data_out_B_for_next2 = Data_Output_B_Mem86;
		
			data_out_A_for_next3 = Data_Output_A_Mem87;
			data_out_B_for_next3 = Data_Output_B_Mem87;
		
			data_out_A_for_next4 = Data_Output_A_Mem88;
			data_out_B_for_next4 = Data_Output_B_Mem88;
		
			data_out_A_for_next5 = Data_Output_A_Mem89;
			data_out_B_for_next5 = Data_Output_B_Mem89;
		
			data_out_A_for_next6 = Data_Output_A_Mem90;
			data_out_B_for_next6 = Data_Output_B_Mem90;
		
			data_out_A_for_next7 = Data_Output_A_Mem91;
			data_out_B_for_next7 = Data_Output_B_Mem91;
		end
		5'd14:
		begin
			data_out_for_previous1 = Data_Output_B_Mem99;
			data_out_for_previous2 = Data_Output_B_Mem100;
			data_out_for_previous3 = Data_Output_B_Mem101;
			data_out_for_previous4 = Data_Output_B_Mem102;
			data_out_for_previous5 = Data_Output_B_Mem103;
			data_out_for_previous6 = Data_Output_B_Mem104;
			data_out_for_previous7 = Data_Output_B_Mem105;
		
			data_out_A_for_next1 = Data_Output_A_Mem92;
			data_out_B_for_next1 = Data_Output_B_Mem92;
		
			data_out_A_for_next2 = Data_Output_A_Mem93;
			data_out_B_for_next2 = Data_Output_B_Mem93;
		
			data_out_A_for_next3 = Data_Output_A_Mem94;
			data_out_B_for_next3 = Data_Output_B_Mem94;
		
			data_out_A_for_next4 = Data_Output_A_Mem95;
			data_out_B_for_next4 = Data_Output_B_Mem95;
		
			data_out_A_for_next5 = Data_Output_A_Mem96;
			data_out_B_for_next5 = Data_Output_B_Mem96;
		
			data_out_A_for_next6 = Data_Output_A_Mem97;
			data_out_B_for_next6 = Data_Output_B_Mem97;
		
			data_out_A_for_next7 = Data_Output_A_Mem98;
			data_out_B_for_next7 = Data_Output_B_Mem98;
		end
		5'd15:
		begin
			data_out_for_previous1 = Data_Output_B_Mem106;
			data_out_for_previous2 = Data_Output_B_Mem107;
			data_out_for_previous3 = Data_Output_B_Mem108;
			data_out_for_previous4 = Data_Output_B_Mem109;
			data_out_for_previous5 = Data_Output_B_Mem110;
			data_out_for_previous6 = Data_Output_B_Mem111;
			data_out_for_previous7 = Data_Output_B_Mem112;
		
			data_out_A_for_next1 = Data_Output_A_Mem99;
			data_out_B_for_next1 = Data_Output_B_Mem99;
		
			data_out_A_for_next2 = Data_Output_A_Mem100;
			data_out_B_for_next2 = Data_Output_B_Mem100;
		
			data_out_A_for_next3 = Data_Output_A_Mem101;
			data_out_B_for_next3 = Data_Output_B_Mem101;
		
			data_out_A_for_next4 = Data_Output_A_Mem102;
			data_out_B_for_next4 = Data_Output_B_Mem102;
		
			data_out_A_for_next5 = Data_Output_A_Mem103;
			data_out_B_for_next5 = Data_Output_B_Mem103;
		
			data_out_A_for_next6 = Data_Output_A_Mem104;
			data_out_B_for_next6 = Data_Output_B_Mem104;
		
			data_out_A_for_next7 = Data_Output_A_Mem105;
			data_out_B_for_next7 = Data_Output_B_Mem105;
		end
		5'd16:
		begin
			data_out_for_previous1 = Data_Output_B_Mem113;
			data_out_for_previous2 = Data_Output_B_Mem114;
			data_out_for_previous3 = Data_Output_B_Mem115;
			data_out_for_previous4 = Data_Output_B_Mem116;
			data_out_for_previous5 = Data_Output_B_Mem117;
			data_out_for_previous6 = Data_Output_B_Mem118;
			data_out_for_previous7 = Data_Output_B_Mem119;
		
			data_out_A_for_next1 = Data_Output_A_Mem106;
			data_out_B_for_next1 = Data_Output_B_Mem106;
		
			data_out_A_for_next2 = Data_Output_A_Mem107;
			data_out_B_for_next2 = Data_Output_B_Mem107;
		
			data_out_A_for_next3 = Data_Output_A_Mem108;
			data_out_B_for_next3 = Data_Output_B_Mem108;
		
			data_out_A_for_next4 = Data_Output_A_Mem109;
			data_out_B_for_next4 = Data_Output_B_Mem109;
		
			data_out_A_for_next5 = Data_Output_A_Mem110;
			data_out_B_for_next5 = Data_Output_B_Mem110;
		
			data_out_A_for_next6 = Data_Output_A_Mem111;
			data_out_B_for_next6 = Data_Output_B_Mem111;
		
			data_out_A_for_next7 = Data_Output_A_Mem112;
			data_out_B_for_next7 = Data_Output_B_Mem112;
		end
		5'd17:
		begin
			data_out_for_previous1 = Data_Output_B_Mem120;
			data_out_for_previous2 = Data_Output_B_Mem121;
			data_out_for_previous3 = Data_Output_B_Mem122;
			data_out_for_previous4 = Data_Output_B_Mem123;
			data_out_for_previous5 = Data_Output_B_Mem124;
			data_out_for_previous6 = Data_Output_B_Mem125;
			data_out_for_previous7 = Data_Output_B_Mem126;
		
			data_out_A_for_next1 = Data_Output_A_Mem113;
			data_out_B_for_next1 = Data_Output_B_Mem113;
		
			data_out_A_for_next2 = Data_Output_A_Mem114;
			data_out_B_for_next2 = Data_Output_B_Mem114;
		
			data_out_A_for_next3 = Data_Output_A_Mem115;
			data_out_B_for_next3 = Data_Output_B_Mem115;
		
			data_out_A_for_next4 = Data_Output_A_Mem116;
			data_out_B_for_next4 = Data_Output_B_Mem116;
		
			data_out_A_for_next5 = Data_Output_A_Mem117;
			data_out_B_for_next5 = Data_Output_B_Mem117;
		
			data_out_A_for_next6 = Data_Output_A_Mem118;
			data_out_B_for_next6 = Data_Output_B_Mem118;
		
			data_out_A_for_next7 = Data_Output_A_Mem119;
			data_out_B_for_next7 = Data_Output_B_Mem119;
		end
		5'd18:
		begin
			data_out_for_previous1 = Data_Output_B_Mem127;
			data_out_for_previous2 = Data_Output_B_Mem128;
			data_out_for_previous3 = Data_Output_B_Mem129;
			data_out_for_previous4 = Data_Output_B_Mem130;
			data_out_for_previous5 = Data_Output_B_Mem131;
			data_out_for_previous6 = Data_Output_B_Mem132;
			data_out_for_previous7 = Data_Output_B_Mem133;
		
			data_out_A_for_next1 = Data_Output_A_Mem120;
			data_out_B_for_next1 = Data_Output_B_Mem120;
		
			data_out_A_for_next2 = Data_Output_A_Mem121;
			data_out_B_for_next2 = Data_Output_B_Mem121;
		
			data_out_A_for_next3 = Data_Output_A_Mem122;
			data_out_B_for_next3 = Data_Output_B_Mem122;
		
			data_out_A_for_next4 = Data_Output_A_Mem123;
			data_out_B_for_next4 = Data_Output_B_Mem123;
		
			data_out_A_for_next5 = Data_Output_A_Mem124;
			data_out_B_for_next5 = Data_Output_B_Mem124;
		
			data_out_A_for_next6 = Data_Output_A_Mem125;
			data_out_B_for_next6 = Data_Output_B_Mem125;
		
			data_out_A_for_next7 = Data_Output_A_Mem126;
			data_out_B_for_next7 = Data_Output_B_Mem126;
		end
		5'd19:
		begin
			data_out_for_previous1 = Data_Output_B_Mem134;
			data_out_for_previous2 = Data_Output_B_Mem135;
			data_out_for_previous3 = Data_Output_B_Mem136;
			data_out_for_previous4 = Data_Output_B_Mem137;
			data_out_for_previous5 = Data_Output_B_Mem138;
			data_out_for_previous6 = Data_Output_B_Mem139;
			data_out_for_previous7 = Data_Output_B_Mem140;
		
			data_out_A_for_next1 = Data_Output_A_Mem127;
			data_out_B_for_next1 = Data_Output_B_Mem127;
		
			data_out_A_for_next2 = Data_Output_A_Mem128;
			data_out_B_for_next2 = Data_Output_B_Mem128;
		
			data_out_A_for_next3 = Data_Output_A_Mem129;
			data_out_B_for_next3 = Data_Output_B_Mem129;
		
			data_out_A_for_next4 = Data_Output_A_Mem130;
			data_out_B_for_next4 = Data_Output_B_Mem130;
		
			data_out_A_for_next5 = Data_Output_A_Mem131;
			data_out_B_for_next5 = Data_Output_B_Mem131;
		
			data_out_A_for_next6 = Data_Output_A_Mem132;
			data_out_B_for_next6 = Data_Output_B_Mem132;
		
			data_out_A_for_next7 = Data_Output_A_Mem133;
			data_out_B_for_next7 = Data_Output_B_Mem133;
		end
		5'd20:
		begin
			data_out_for_previous1 = Data_Output_B_Mem141;
			data_out_for_previous2 = Data_Output_B_Mem142;
			data_out_for_previous3 = Data_Output_B_Mem143;
			data_out_for_previous4 = Data_Output_B_Mem144;
			data_out_for_previous5 = Data_Output_B_Mem145;
			data_out_for_previous6 = Data_Output_B_Mem146;
			data_out_for_previous7 = Data_Output_B_Mem147;
		
			data_out_A_for_next1 = Data_Output_A_Mem134;
			data_out_B_for_next1 = Data_Output_B_Mem134;
		
			data_out_A_for_next2 = Data_Output_A_Mem135;
			data_out_B_for_next2 = Data_Output_B_Mem135;
		
			data_out_A_for_next3 = Data_Output_A_Mem136;
			data_out_B_for_next3 = Data_Output_B_Mem136;
		
			data_out_A_for_next4 = Data_Output_A_Mem137;
			data_out_B_for_next4 = Data_Output_B_Mem137;
		
			data_out_A_for_next5 = Data_Output_A_Mem138;
			data_out_B_for_next5 = Data_Output_B_Mem138;
		
			data_out_A_for_next6 = Data_Output_A_Mem139;
			data_out_B_for_next6 = Data_Output_B_Mem139;
		
			data_out_A_for_next7 = Data_Output_A_Mem140;
			data_out_B_for_next7 = Data_Output_B_Mem140;
		end
		5'd21:
		begin
			data_out_for_previous1 = Data_Output_B_Mem148;
			data_out_for_previous2 = Data_Output_B_Mem149;
			data_out_for_previous3 = Data_Output_B_Mem150;
			data_out_for_previous4 = Data_Output_B_Mem151;
			data_out_for_previous5 = Data_Output_B_Mem152;
			data_out_for_previous6 = Data_Output_B_Mem153;
			data_out_for_previous7 = Data_Output_B_Mem154;
		
			data_out_A_for_next1 = Data_Output_A_Mem141;
			data_out_B_for_next1 = Data_Output_B_Mem141;
		
			data_out_A_for_next2 = Data_Output_A_Mem142;
			data_out_B_for_next2 = Data_Output_B_Mem142;
		
			data_out_A_for_next3 = Data_Output_A_Mem143;
			data_out_B_for_next3 = Data_Output_B_Mem143;
		
			data_out_A_for_next4 = Data_Output_A_Mem144;
			data_out_B_for_next4 = Data_Output_B_Mem144;
		
			data_out_A_for_next5 = Data_Output_A_Mem145;
			data_out_B_for_next5 = Data_Output_B_Mem145;
		
			data_out_A_for_next6 = Data_Output_A_Mem146;
			data_out_B_for_next6 = Data_Output_B_Mem146;
		
			data_out_A_for_next7 = Data_Output_A_Mem147;
			data_out_B_for_next7 = Data_Output_B_Mem147;
		end
		5'd22:
		begin
			data_out_for_previous1 = Data_Output_B_Mem155;
			data_out_for_previous2 = Data_Output_B_Mem156;
			data_out_for_previous3 = Data_Output_B_Mem157;
			data_out_for_previous4 = Data_Output_B_Mem158;
			data_out_for_previous5 = Data_Output_B_Mem159;
			data_out_for_previous6 = Data_Output_B_Mem160;
			data_out_for_previous7 = Data_Output_B_Mem161;
		
			data_out_A_for_next1 = Data_Output_A_Mem148;
			data_out_B_for_next1 = Data_Output_B_Mem148;
		
			data_out_A_for_next2 = Data_Output_A_Mem149;
			data_out_B_for_next2 = Data_Output_B_Mem149;
		
			data_out_A_for_next3 = Data_Output_A_Mem150;
			data_out_B_for_next3 = Data_Output_B_Mem150;
		
			data_out_A_for_next4 = Data_Output_A_Mem151;
			data_out_B_for_next4 = Data_Output_B_Mem151;
		
			data_out_A_for_next5 = Data_Output_A_Mem152;
			data_out_B_for_next5 = Data_Output_B_Mem152;
		
			data_out_A_for_next6 = Data_Output_A_Mem153;
			data_out_B_for_next6 = Data_Output_B_Mem153;
		
			data_out_A_for_next7 = Data_Output_A_Mem154;
			data_out_B_for_next7 = Data_Output_B_Mem154;
		end
		5'd23:
		begin
			data_out_for_previous1 = Data_Output_B_Mem162;
			data_out_for_previous2 = Data_Output_B_Mem163;
			data_out_for_previous3 = Data_Output_B_Mem164;
			data_out_for_previous4 = Data_Output_B_Mem165;
			data_out_for_previous5 = Data_Output_B_Mem166;
			data_out_for_previous6 = Data_Output_B_Mem167;
			data_out_for_previous7 = Data_Output_B_Mem168;
		
			data_out_A_for_next1 = Data_Output_A_Mem155;
			data_out_B_for_next1 = Data_Output_B_Mem155;
		
			data_out_A_for_next2 = Data_Output_A_Mem156;
			data_out_B_for_next2 = Data_Output_B_Mem156;
		
			data_out_A_for_next3 = Data_Output_A_Mem157;
			data_out_B_for_next3 = Data_Output_B_Mem157;
		
			data_out_A_for_next4 = Data_Output_A_Mem158;
			data_out_B_for_next4 = Data_Output_B_Mem158;
		
			data_out_A_for_next5 = Data_Output_A_Mem159;
			data_out_B_for_next5 = Data_Output_B_Mem159;
		
			data_out_A_for_next6 = Data_Output_A_Mem160;
			data_out_B_for_next6 = Data_Output_B_Mem160;
		
			data_out_A_for_next7 = Data_Output_A_Mem161;
			data_out_B_for_next7 = Data_Output_B_Mem161;
		end
		5'd24:
		begin
			data_out_for_previous1 = Data_Output_B_Mem169;
			data_out_for_previous2 = Data_Output_B_Mem170;
			data_out_for_previous3 = Data_Output_B_Mem171;
			data_out_for_previous4 = Data_Output_B_Mem172;
			data_out_for_previous5 = Data_Output_B_Mem173;
			data_out_for_previous6 = Data_Output_B_Mem174;
			data_out_for_previous7 = Data_Output_B_Mem175;
		
			data_out_A_for_next1 = Data_Output_A_Mem162;
			data_out_B_for_next1 = Data_Output_B_Mem162;
		
			data_out_A_for_next2 = Data_Output_A_Mem163;
			data_out_B_for_next2 = Data_Output_B_Mem163;
		
			data_out_A_for_next3 = Data_Output_A_Mem164;
			data_out_B_for_next3 = Data_Output_B_Mem164;
		
			data_out_A_for_next4 = Data_Output_A_Mem165;
			data_out_B_for_next4 = Data_Output_B_Mem165;
		
			data_out_A_for_next5 = Data_Output_A_Mem166;
			data_out_B_for_next5 = Data_Output_B_Mem166;
		
			data_out_A_for_next6 = Data_Output_A_Mem167;
			data_out_B_for_next6 = Data_Output_B_Mem167;
		
			data_out_A_for_next7 = Data_Output_A_Mem168;
			data_out_B_for_next7 = Data_Output_B_Mem168;
		end
		5'd25:
		begin
			data_out_for_previous1 = Data_Output_B_Mem176;
			data_out_for_previous2 = Data_Output_B_Mem177;
			data_out_for_previous3 = Data_Output_B_Mem178;
			data_out_for_previous4 = Data_Output_B_Mem179;
			data_out_for_previous5 = Data_Output_B_Mem180;
			data_out_for_previous6 = Data_Output_B_Mem181;
			data_out_for_previous7 = Data_Output_B_Mem182;
		
			data_out_A_for_next1 = Data_Output_A_Mem169;
			data_out_B_for_next1 = Data_Output_B_Mem169;
		
			data_out_A_for_next2 = Data_Output_A_Mem170;
			data_out_B_for_next2 = Data_Output_B_Mem170;
		
			data_out_A_for_next3 = Data_Output_A_Mem171;
			data_out_B_for_next3 = Data_Output_B_Mem171;
		
			data_out_A_for_next4 = Data_Output_A_Mem172;
			data_out_B_for_next4 = Data_Output_B_Mem172;
		
			data_out_A_for_next5 = Data_Output_A_Mem173;
			data_out_B_for_next5 = Data_Output_B_Mem173;
		
			data_out_A_for_next6 = Data_Output_A_Mem174;
			data_out_B_for_next6 = Data_Output_B_Mem174;
		
			data_out_A_for_next7 = Data_Output_A_Mem175;
			data_out_B_for_next7 = Data_Output_B_Mem175;
		end
		5'd26:
		begin
			data_out_for_previous1 = Data_Output_B_Mem183;
			data_out_for_previous2 = Data_Output_B_Mem184;
			data_out_for_previous3 = Data_Output_B_Mem185;
			data_out_for_previous4 = Data_Output_B_Mem186;
			data_out_for_previous5 = Data_Output_B_Mem187;
			data_out_for_previous6 = Data_Output_B_Mem188;
			data_out_for_previous7 = Data_Output_B_Mem189;
		
			data_out_A_for_next1 = Data_Output_A_Mem176;
			data_out_B_for_next1 = Data_Output_B_Mem176;
		
			data_out_A_for_next2 = Data_Output_A_Mem177;
			data_out_B_for_next2 = Data_Output_B_Mem177;
		
			data_out_A_for_next3 = Data_Output_A_Mem178;
			data_out_B_for_next3 = Data_Output_B_Mem178;
		
			data_out_A_for_next4 = Data_Output_A_Mem179;
			data_out_B_for_next4 = Data_Output_B_Mem179;
		
			data_out_A_for_next5 = Data_Output_A_Mem180;
			data_out_B_for_next5 = Data_Output_B_Mem180;
		
			data_out_A_for_next6 = Data_Output_A_Mem181;
			data_out_B_for_next6 = Data_Output_B_Mem181;
		
			data_out_A_for_next7 = Data_Output_A_Mem182;
			data_out_B_for_next7 = Data_Output_B_Mem182;
		end
		5'd27:
		begin
			data_out_for_previous1 = Data_Output_B_Mem190;
			data_out_for_previous2 = Data_Output_B_Mem191;
			data_out_for_previous3 = Data_Output_B_Mem192;
			data_out_for_previous4 = Data_Output_B_Mem193;
			data_out_for_previous5 = Data_Output_B_Mem194;
			data_out_for_previous6 = Data_Output_B_Mem195;
			data_out_for_previous7 = Data_Output_B_Mem196;
		
			data_out_A_for_next1 = Data_Output_A_Mem183;
			data_out_B_for_next1 = Data_Output_B_Mem183;
		
			data_out_A_for_next2 = Data_Output_A_Mem184;
			data_out_B_for_next2 = Data_Output_B_Mem184;
		
			data_out_A_for_next3 = Data_Output_A_Mem185;
			data_out_B_for_next3 = Data_Output_B_Mem185;
		
			data_out_A_for_next4 = Data_Output_A_Mem186;
			data_out_B_for_next4 = Data_Output_B_Mem186;
		
			data_out_A_for_next5 = Data_Output_A_Mem187;
			data_out_B_for_next5 = Data_Output_B_Mem187;
		
			data_out_A_for_next6 = Data_Output_A_Mem188;
			data_out_B_for_next6 = Data_Output_B_Mem188;
		
			data_out_A_for_next7 = Data_Output_A_Mem189;
			data_out_B_for_next7 = Data_Output_B_Mem189;
		end
		default:
		begin
			data_out_for_previous1 = Data_Output_B_Mem197;
			data_out_for_previous2 = Data_Output_B_Mem198;
			data_out_for_previous3 = Data_Output_B_Mem199;
			data_out_for_previous4 = Data_Output_B_Mem200;
			data_out_for_previous5 = 0;
			data_out_for_previous6 = 0;
			data_out_for_previous7 = 0;
		
			data_out_A_for_next1 = Data_Output_A_Mem190;
			data_out_B_for_next1 = Data_Output_B_Mem190;
		
			data_out_A_for_next2 = Data_Output_A_Mem191;
			data_out_B_for_next2 = Data_Output_B_Mem191;
		
			data_out_A_for_next3 = Data_Output_A_Mem192;
			data_out_B_for_next3 = Data_Output_B_Mem192;
		
			data_out_A_for_next4 = Data_Output_A_Mem193;
			data_out_B_for_next4 = Data_Output_B_Mem193;
		
			data_out_A_for_next5 = Data_Output_A_Mem194;
			data_out_B_for_next5 = Data_Output_B_Mem194;
		
			data_out_A_for_next6 = Data_Output_A_Mem195;
			data_out_B_for_next6 = Data_Output_B_Mem195;
		
			data_out_A_for_next7 = Data_Output_A_Mem196;
			data_out_B_for_next7 = Data_Output_B_Mem196;
		end
		
		endcase
		
	end
	
mem_unit #( .DATA_WIDTH(DATA_WIDTH),.IFM_SIZE(IFM_SIZE))
M1(  .clk(clk),
      .Data_Input_A_Mem1 (data_in_from_previous1),
      .Data_Input_B_Mem1 ('b0),
      .Data_Input_A_Mem2 (data_in_from_previous2),
      .Data_Input_B_Mem2 ('b0),
      .Data_Input_A_Mem3 (data_in_from_previous3),
      .Data_Input_B_Mem3 ('b0),
      .Data_Input_A_Mem4 (data_in_from_previous4),
      .Data_Input_B_Mem4 ('b0),
      .Data_Input_A_Mem5 (data_in_from_previous5),
      .Data_Input_B_Mem5 ('b0),
      .Data_Input_A_Mem6 (data_in_from_previous6),
      .Data_Input_B_Mem6 ('b0),
      .Data_Input_A_Mem7 (data_in_from_previous7),
      .Data_Input_B_Mem7 ('b0),
	
      .Address_A ( ifm_address_write_previous_dMuxOut1 | ifm_address_read_A_next_dMuxOut2 ),
      .Address_B ( ifm_address_read_previous_dMuxOut1  | ifm_address_read_B_next_dMuxOut2 ),  
	
      .Enable_Write_A_Mem (ifm_enable_write_previous_dMuxOut1),
      .Enable_Read_A_Mem  (ifm_enable_read_A_next_dMuxOut2),
      .Enable_Write_B_Mem (1'b0),
      .Enable_Read_B_Mem  (ifm_enable_read_previous_dMuxOut1 | ifm_enable_read_B_next_dMuxOut2),
	  
      .Data_Output_A_Mem1 (Data_Output_A_Mem1),
      .Data_Output_B_Mem1 (Data_Output_B_Mem1),
      .Data_Output_A_Mem2 (Data_Output_A_Mem2),
      .Data_Output_B_Mem2 (Data_Output_B_Mem2),
      .Data_Output_A_Mem3 (Data_Output_A_Mem3),
      .Data_Output_B_Mem3 (Data_Output_B_Mem3),
      .Data_Output_A_Mem4 (Data_Output_A_Mem4),
      .Data_Output_B_Mem4 (Data_Output_B_Mem4),
      .Data_Output_A_Mem5 (Data_Output_A_Mem5),
      .Data_Output_B_Mem5 (Data_Output_B_Mem5),
      .Data_Output_A_Mem6 (Data_Output_A_Mem6),
      .Data_Output_B_Mem6 (Data_Output_B_Mem6),
      .Data_Output_A_Mem7 (Data_Output_A_Mem7),
      .Data_Output_B_Mem7 (Data_Output_B_Mem7)
	  );
	
mem_unit #( .DATA_WIDTH(DATA_WIDTH),.IFM_SIZE(IFM_SIZE))
M2(  .clk(clk),
      .Data_Input_A_Mem1 (data_in_from_previous1),
      .Data_Input_B_Mem1 ('b0),
      .Data_Input_A_Mem2 (data_in_from_previous2),
      .Data_Input_B_Mem2 ('b0),
      .Data_Input_A_Mem3 (data_in_from_previous3),
      .Data_Input_B_Mem3 ('b0),
      .Data_Input_A_Mem4 (data_in_from_previous4),
      .Data_Input_B_Mem4 ('b0),
      .Data_Input_A_Mem5 (data_in_from_previous5),
      .Data_Input_B_Mem5 ('b0),
      .Data_Input_A_Mem6 (data_in_from_previous6),
      .Data_Input_B_Mem6 ('b0),
      .Data_Input_A_Mem7 (data_in_from_previous7),
      .Data_Input_B_Mem7 ('b0),
	
      .Address_A ( ifm_address_write_previous_dMuxOut2 | ifm_address_read_A_next_dMuxOut3 ),
      .Address_B ( ifm_address_read_previous_dMuxOut2  | ifm_address_read_B_next_dMuxOut3 ),  
	
      .Enable_Write_A_Mem (ifm_enable_write_previous_dMuxOut2),
      .Enable_Read_A_Mem  (ifm_enable_read_A_next_dMuxOut3),
      .Enable_Write_B_Mem (1'b0),
      .Enable_Read_B_Mem  (ifm_enable_read_previous_dMuxOut2 | ifm_enable_read_B_next_dMuxOut3),
	  
      .Data_Output_A_Mem1 (Data_Output_A_Mem8),
      .Data_Output_B_Mem1 (Data_Output_B_Mem8),
      .Data_Output_A_Mem2 (Data_Output_A_Mem9),
      .Data_Output_B_Mem2 (Data_Output_B_Mem9),
      .Data_Output_A_Mem3 (Data_Output_A_Mem10),
      .Data_Output_B_Mem3 (Data_Output_B_Mem10),
      .Data_Output_A_Mem4 (Data_Output_A_Mem11),
      .Data_Output_B_Mem4 (Data_Output_B_Mem11),
      .Data_Output_A_Mem5 (Data_Output_A_Mem12),
      .Data_Output_B_Mem5 (Data_Output_B_Mem12),
      .Data_Output_A_Mem6 (Data_Output_A_Mem13),
      .Data_Output_B_Mem6 (Data_Output_B_Mem13),
      .Data_Output_A_Mem7 (Data_Output_A_Mem14),
      .Data_Output_B_Mem7 (Data_Output_B_Mem14)
	  );
	
mem_unit #( .DATA_WIDTH(DATA_WIDTH),.IFM_SIZE(IFM_SIZE))
M3(  .clk(clk),
      .Data_Input_A_Mem1 (data_in_from_previous1),
      .Data_Input_B_Mem1 ('b0),
      .Data_Input_A_Mem2 (data_in_from_previous2),
      .Data_Input_B_Mem2 ('b0),
      .Data_Input_A_Mem3 (data_in_from_previous3),
      .Data_Input_B_Mem3 ('b0),
      .Data_Input_A_Mem4 (data_in_from_previous4),
      .Data_Input_B_Mem4 ('b0),
      .Data_Input_A_Mem5 (data_in_from_previous5),
      .Data_Input_B_Mem5 ('b0),
      .Data_Input_A_Mem6 (data_in_from_previous6),
      .Data_Input_B_Mem6 ('b0),
      .Data_Input_A_Mem7 (data_in_from_previous7),
      .Data_Input_B_Mem7 ('b0),
	
      .Address_A ( ifm_address_write_previous_dMuxOut3 | ifm_address_read_A_next_dMuxOut4 ),
      .Address_B ( ifm_address_read_previous_dMuxOut3  | ifm_address_read_B_next_dMuxOut4 ),  
	
      .Enable_Write_A_Mem (ifm_enable_write_previous_dMuxOut3),
      .Enable_Read_A_Mem  (ifm_enable_read_A_next_dMuxOut4),
      .Enable_Write_B_Mem (1'b0),
      .Enable_Read_B_Mem  (ifm_enable_read_previous_dMuxOut3 | ifm_enable_read_B_next_dMuxOut4),
	  
      .Data_Output_A_Mem1 (Data_Output_A_Mem15),
      .Data_Output_B_Mem1 (Data_Output_B_Mem15),
      .Data_Output_A_Mem2 (Data_Output_A_Mem16),
      .Data_Output_B_Mem2 (Data_Output_B_Mem16),
      .Data_Output_A_Mem3 (Data_Output_A_Mem17),
      .Data_Output_B_Mem3 (Data_Output_B_Mem17),
      .Data_Output_A_Mem4 (Data_Output_A_Mem18),
      .Data_Output_B_Mem4 (Data_Output_B_Mem18),
      .Data_Output_A_Mem5 (Data_Output_A_Mem19),
      .Data_Output_B_Mem5 (Data_Output_B_Mem19),
      .Data_Output_A_Mem6 (Data_Output_A_Mem20),
      .Data_Output_B_Mem6 (Data_Output_B_Mem20),
      .Data_Output_A_Mem7 (Data_Output_A_Mem21),
      .Data_Output_B_Mem7 (Data_Output_B_Mem21)
	  );
	
mem_unit #( .DATA_WIDTH(DATA_WIDTH),.IFM_SIZE(IFM_SIZE))
M4(  .clk(clk),
      .Data_Input_A_Mem1 (data_in_from_previous1),
      .Data_Input_B_Mem1 ('b0),
      .Data_Input_A_Mem2 (data_in_from_previous2),
      .Data_Input_B_Mem2 ('b0),
      .Data_Input_A_Mem3 (data_in_from_previous3),
      .Data_Input_B_Mem3 ('b0),
      .Data_Input_A_Mem4 (data_in_from_previous4),
      .Data_Input_B_Mem4 ('b0),
      .Data_Input_A_Mem5 (data_in_from_previous5),
      .Data_Input_B_Mem5 ('b0),
      .Data_Input_A_Mem6 (data_in_from_previous6),
      .Data_Input_B_Mem6 ('b0),
      .Data_Input_A_Mem7 (data_in_from_previous7),
      .Data_Input_B_Mem7 ('b0),
	
      .Address_A ( ifm_address_write_previous_dMuxOut4 | ifm_address_read_A_next_dMuxOut5 ),
      .Address_B ( ifm_address_read_previous_dMuxOut4  | ifm_address_read_B_next_dMuxOut5 ),  
	
      .Enable_Write_A_Mem (ifm_enable_write_previous_dMuxOut4),
      .Enable_Read_A_Mem  (ifm_enable_read_A_next_dMuxOut5),
      .Enable_Write_B_Mem (1'b0),
      .Enable_Read_B_Mem  (ifm_enable_read_previous_dMuxOut4 | ifm_enable_read_B_next_dMuxOut5),
	  
      .Data_Output_A_Mem1 (Data_Output_A_Mem22),
      .Data_Output_B_Mem1 (Data_Output_B_Mem22),
      .Data_Output_A_Mem2 (Data_Output_A_Mem23),
      .Data_Output_B_Mem2 (Data_Output_B_Mem23),
      .Data_Output_A_Mem3 (Data_Output_A_Mem24),
      .Data_Output_B_Mem3 (Data_Output_B_Mem24),
      .Data_Output_A_Mem4 (Data_Output_A_Mem25),
      .Data_Output_B_Mem4 (Data_Output_B_Mem25),
      .Data_Output_A_Mem5 (Data_Output_A_Mem26),
      .Data_Output_B_Mem5 (Data_Output_B_Mem26),
      .Data_Output_A_Mem6 (Data_Output_A_Mem27),
      .Data_Output_B_Mem6 (Data_Output_B_Mem27),
      .Data_Output_A_Mem7 (Data_Output_A_Mem28),
      .Data_Output_B_Mem7 (Data_Output_B_Mem28)
	  );
	
mem_unit #( .DATA_WIDTH(DATA_WIDTH),.IFM_SIZE(IFM_SIZE))
M5(  .clk(clk),
      .Data_Input_A_Mem1 (data_in_from_previous1),
      .Data_Input_B_Mem1 ('b0),
      .Data_Input_A_Mem2 (data_in_from_previous2),
      .Data_Input_B_Mem2 ('b0),
      .Data_Input_A_Mem3 (data_in_from_previous3),
      .Data_Input_B_Mem3 ('b0),
      .Data_Input_A_Mem4 (data_in_from_previous4),
      .Data_Input_B_Mem4 ('b0),
      .Data_Input_A_Mem5 (data_in_from_previous5),
      .Data_Input_B_Mem5 ('b0),
      .Data_Input_A_Mem6 (data_in_from_previous6),
      .Data_Input_B_Mem6 ('b0),
      .Data_Input_A_Mem7 (data_in_from_previous7),
      .Data_Input_B_Mem7 ('b0),
	
      .Address_A ( ifm_address_write_previous_dMuxOut5 | ifm_address_read_A_next_dMuxOut6 ),
      .Address_B ( ifm_address_read_previous_dMuxOut5  | ifm_address_read_B_next_dMuxOut6 ),  
	
      .Enable_Write_A_Mem (ifm_enable_write_previous_dMuxOut5),
      .Enable_Read_A_Mem  (ifm_enable_read_A_next_dMuxOut6),
      .Enable_Write_B_Mem (1'b0),
      .Enable_Read_B_Mem  (ifm_enable_read_previous_dMuxOut5 | ifm_enable_read_B_next_dMuxOut6),
	  
      .Data_Output_A_Mem1 (Data_Output_A_Mem29),
      .Data_Output_B_Mem1 (Data_Output_B_Mem29),
      .Data_Output_A_Mem2 (Data_Output_A_Mem30),
      .Data_Output_B_Mem2 (Data_Output_B_Mem30),
      .Data_Output_A_Mem3 (Data_Output_A_Mem31),
      .Data_Output_B_Mem3 (Data_Output_B_Mem31),
      .Data_Output_A_Mem4 (Data_Output_A_Mem32),
      .Data_Output_B_Mem4 (Data_Output_B_Mem32),
      .Data_Output_A_Mem5 (Data_Output_A_Mem33),
      .Data_Output_B_Mem5 (Data_Output_B_Mem33),
      .Data_Output_A_Mem6 (Data_Output_A_Mem34),
      .Data_Output_B_Mem6 (Data_Output_B_Mem34),
      .Data_Output_A_Mem7 (Data_Output_A_Mem35),
      .Data_Output_B_Mem7 (Data_Output_B_Mem35)
	  );
	
mem_unit #( .DATA_WIDTH(DATA_WIDTH),.IFM_SIZE(IFM_SIZE))
M6(  .clk(clk),
      .Data_Input_A_Mem1 (data_in_from_previous1),
      .Data_Input_B_Mem1 ('b0),
      .Data_Input_A_Mem2 (data_in_from_previous2),
      .Data_Input_B_Mem2 ('b0),
      .Data_Input_A_Mem3 (data_in_from_previous3),
      .Data_Input_B_Mem3 ('b0),
      .Data_Input_A_Mem4 (data_in_from_previous4),
      .Data_Input_B_Mem4 ('b0),
      .Data_Input_A_Mem5 (data_in_from_previous5),
      .Data_Input_B_Mem5 ('b0),
      .Data_Input_A_Mem6 (data_in_from_previous6),
      .Data_Input_B_Mem6 ('b0),
      .Data_Input_A_Mem7 (data_in_from_previous7),
      .Data_Input_B_Mem7 ('b0),
	
      .Address_A ( ifm_address_write_previous_dMuxOut6 | ifm_address_read_A_next_dMuxOut7 ),
      .Address_B ( ifm_address_read_previous_dMuxOut6  | ifm_address_read_B_next_dMuxOut7 ),  
	
      .Enable_Write_A_Mem (ifm_enable_write_previous_dMuxOut6),
      .Enable_Read_A_Mem  (ifm_enable_read_A_next_dMuxOut7),
      .Enable_Write_B_Mem (1'b0),
      .Enable_Read_B_Mem  (ifm_enable_read_previous_dMuxOut6 | ifm_enable_read_B_next_dMuxOut7),
	  
      .Data_Output_A_Mem1 (Data_Output_A_Mem36),
      .Data_Output_B_Mem1 (Data_Output_B_Mem36),
      .Data_Output_A_Mem2 (Data_Output_A_Mem37),
      .Data_Output_B_Mem2 (Data_Output_B_Mem37),
      .Data_Output_A_Mem3 (Data_Output_A_Mem38),
      .Data_Output_B_Mem3 (Data_Output_B_Mem38),
      .Data_Output_A_Mem4 (Data_Output_A_Mem39),
      .Data_Output_B_Mem4 (Data_Output_B_Mem39),
      .Data_Output_A_Mem5 (Data_Output_A_Mem40),
      .Data_Output_B_Mem5 (Data_Output_B_Mem40),
      .Data_Output_A_Mem6 (Data_Output_A_Mem41),
      .Data_Output_B_Mem6 (Data_Output_B_Mem41),
      .Data_Output_A_Mem7 (Data_Output_A_Mem42),
      .Data_Output_B_Mem7 (Data_Output_B_Mem42)
	  );
	
mem_unit #( .DATA_WIDTH(DATA_WIDTH),.IFM_SIZE(IFM_SIZE))
M7(  .clk(clk),
      .Data_Input_A_Mem1 (data_in_from_previous1),
      .Data_Input_B_Mem1 ('b0),
      .Data_Input_A_Mem2 (data_in_from_previous2),
      .Data_Input_B_Mem2 ('b0),
      .Data_Input_A_Mem3 (data_in_from_previous3),
      .Data_Input_B_Mem3 ('b0),
      .Data_Input_A_Mem4 (data_in_from_previous4),
      .Data_Input_B_Mem4 ('b0),
      .Data_Input_A_Mem5 (data_in_from_previous5),
      .Data_Input_B_Mem5 ('b0),
      .Data_Input_A_Mem6 (data_in_from_previous6),
      .Data_Input_B_Mem6 ('b0),
      .Data_Input_A_Mem7 (data_in_from_previous7),
      .Data_Input_B_Mem7 ('b0),
	
      .Address_A ( ifm_address_write_previous_dMuxOut7 | ifm_address_read_A_next_dMuxOut8 ),
      .Address_B ( ifm_address_read_previous_dMuxOut7  | ifm_address_read_B_next_dMuxOut8 ),  
	
      .Enable_Write_A_Mem (ifm_enable_write_previous_dMuxOut7),
      .Enable_Read_A_Mem  (ifm_enable_read_A_next_dMuxOut8),
      .Enable_Write_B_Mem (1'b0),
      .Enable_Read_B_Mem  (ifm_enable_read_previous_dMuxOut7 | ifm_enable_read_B_next_dMuxOut8),
	  
      .Data_Output_A_Mem1 (Data_Output_A_Mem43),
      .Data_Output_B_Mem1 (Data_Output_B_Mem43),
      .Data_Output_A_Mem2 (Data_Output_A_Mem44),
      .Data_Output_B_Mem2 (Data_Output_B_Mem44),
      .Data_Output_A_Mem3 (Data_Output_A_Mem45),
      .Data_Output_B_Mem3 (Data_Output_B_Mem45),
      .Data_Output_A_Mem4 (Data_Output_A_Mem46),
      .Data_Output_B_Mem4 (Data_Output_B_Mem46),
      .Data_Output_A_Mem5 (Data_Output_A_Mem47),
      .Data_Output_B_Mem5 (Data_Output_B_Mem47),
      .Data_Output_A_Mem6 (Data_Output_A_Mem48),
      .Data_Output_B_Mem6 (Data_Output_B_Mem48),
      .Data_Output_A_Mem7 (Data_Output_A_Mem49),
      .Data_Output_B_Mem7 (Data_Output_B_Mem49)
	  );
	
mem_unit #( .DATA_WIDTH(DATA_WIDTH),.IFM_SIZE(IFM_SIZE))
M8(  .clk(clk),
      .Data_Input_A_Mem1 (data_in_from_previous1),
      .Data_Input_B_Mem1 ('b0),
      .Data_Input_A_Mem2 (data_in_from_previous2),
      .Data_Input_B_Mem2 ('b0),
      .Data_Input_A_Mem3 (data_in_from_previous3),
      .Data_Input_B_Mem3 ('b0),
      .Data_Input_A_Mem4 (data_in_from_previous4),
      .Data_Input_B_Mem4 ('b0),
      .Data_Input_A_Mem5 (data_in_from_previous5),
      .Data_Input_B_Mem5 ('b0),
      .Data_Input_A_Mem6 (data_in_from_previous6),
      .Data_Input_B_Mem6 ('b0),
      .Data_Input_A_Mem7 (data_in_from_previous7),
      .Data_Input_B_Mem7 ('b0),
	
      .Address_A ( ifm_address_write_previous_dMuxOut8 | ifm_address_read_A_next_dMuxOut9 ),
      .Address_B ( ifm_address_read_previous_dMuxOut8  | ifm_address_read_B_next_dMuxOut9 ),  
	
      .Enable_Write_A_Mem (ifm_enable_write_previous_dMuxOut8),
      .Enable_Read_A_Mem  (ifm_enable_read_A_next_dMuxOut9),
      .Enable_Write_B_Mem (1'b0),
      .Enable_Read_B_Mem  (ifm_enable_read_previous_dMuxOut8 | ifm_enable_read_B_next_dMuxOut9),
	  
      .Data_Output_A_Mem1 (Data_Output_A_Mem50),
      .Data_Output_B_Mem1 (Data_Output_B_Mem50),
      .Data_Output_A_Mem2 (Data_Output_A_Mem51),
      .Data_Output_B_Mem2 (Data_Output_B_Mem51),
      .Data_Output_A_Mem3 (Data_Output_A_Mem52),
      .Data_Output_B_Mem3 (Data_Output_B_Mem52),
      .Data_Output_A_Mem4 (Data_Output_A_Mem53),
      .Data_Output_B_Mem4 (Data_Output_B_Mem53),
      .Data_Output_A_Mem5 (Data_Output_A_Mem54),
      .Data_Output_B_Mem5 (Data_Output_B_Mem54),
      .Data_Output_A_Mem6 (Data_Output_A_Mem55),
      .Data_Output_B_Mem6 (Data_Output_B_Mem55),
      .Data_Output_A_Mem7 (Data_Output_A_Mem56),
      .Data_Output_B_Mem7 (Data_Output_B_Mem56)
	  );
	
mem_unit #( .DATA_WIDTH(DATA_WIDTH),.IFM_SIZE(IFM_SIZE))
M9(  .clk(clk),
      .Data_Input_A_Mem1 (data_in_from_previous1),
      .Data_Input_B_Mem1 ('b0),
      .Data_Input_A_Mem2 (data_in_from_previous2),
      .Data_Input_B_Mem2 ('b0),
      .Data_Input_A_Mem3 (data_in_from_previous3),
      .Data_Input_B_Mem3 ('b0),
      .Data_Input_A_Mem4 (data_in_from_previous4),
      .Data_Input_B_Mem4 ('b0),
      .Data_Input_A_Mem5 (data_in_from_previous5),
      .Data_Input_B_Mem5 ('b0),
      .Data_Input_A_Mem6 (data_in_from_previous6),
      .Data_Input_B_Mem6 ('b0),
      .Data_Input_A_Mem7 (data_in_from_previous7),
      .Data_Input_B_Mem7 ('b0),
	
      .Address_A ( ifm_address_write_previous_dMuxOut9 | ifm_address_read_A_next_dMuxOut10 ),
      .Address_B ( ifm_address_read_previous_dMuxOut9  | ifm_address_read_B_next_dMuxOut10 ),  
	
      .Enable_Write_A_Mem (ifm_enable_write_previous_dMuxOut9),
      .Enable_Read_A_Mem  (ifm_enable_read_A_next_dMuxOut10),
      .Enable_Write_B_Mem (1'b0),
      .Enable_Read_B_Mem  (ifm_enable_read_previous_dMuxOut9 | ifm_enable_read_B_next_dMuxOut10),
	  
      .Data_Output_A_Mem1 (Data_Output_A_Mem57),
      .Data_Output_B_Mem1 (Data_Output_B_Mem57),
      .Data_Output_A_Mem2 (Data_Output_A_Mem58),
      .Data_Output_B_Mem2 (Data_Output_B_Mem58),
      .Data_Output_A_Mem3 (Data_Output_A_Mem59),
      .Data_Output_B_Mem3 (Data_Output_B_Mem59),
      .Data_Output_A_Mem4 (Data_Output_A_Mem60),
      .Data_Output_B_Mem4 (Data_Output_B_Mem60),
      .Data_Output_A_Mem5 (Data_Output_A_Mem61),
      .Data_Output_B_Mem5 (Data_Output_B_Mem61),
      .Data_Output_A_Mem6 (Data_Output_A_Mem62),
      .Data_Output_B_Mem6 (Data_Output_B_Mem62),
      .Data_Output_A_Mem7 (Data_Output_A_Mem63),
      .Data_Output_B_Mem7 (Data_Output_B_Mem63)
	  );
	
mem_unit #( .DATA_WIDTH(DATA_WIDTH),.IFM_SIZE(IFM_SIZE))
M10(  .clk(clk),
      .Data_Input_A_Mem1 (data_in_from_previous1),
      .Data_Input_B_Mem1 ('b0),
      .Data_Input_A_Mem2 (data_in_from_previous2),
      .Data_Input_B_Mem2 ('b0),
      .Data_Input_A_Mem3 (data_in_from_previous3),
      .Data_Input_B_Mem3 ('b0),
      .Data_Input_A_Mem4 (data_in_from_previous4),
      .Data_Input_B_Mem4 ('b0),
      .Data_Input_A_Mem5 (data_in_from_previous5),
      .Data_Input_B_Mem5 ('b0),
      .Data_Input_A_Mem6 (data_in_from_previous6),
      .Data_Input_B_Mem6 ('b0),
      .Data_Input_A_Mem7 (data_in_from_previous7),
      .Data_Input_B_Mem7 ('b0),
	
      .Address_A ( ifm_address_write_previous_dMuxOut10 | ifm_address_read_A_next_dMuxOut11 ),
      .Address_B ( ifm_address_read_previous_dMuxOut10  | ifm_address_read_B_next_dMuxOut11 ),  
	
      .Enable_Write_A_Mem (ifm_enable_write_previous_dMuxOut10),
      .Enable_Read_A_Mem  (ifm_enable_read_A_next_dMuxOut11),
      .Enable_Write_B_Mem (1'b0),
      .Enable_Read_B_Mem  (ifm_enable_read_previous_dMuxOut10 | ifm_enable_read_B_next_dMuxOut11),
	  
      .Data_Output_A_Mem1 (Data_Output_A_Mem64),
      .Data_Output_B_Mem1 (Data_Output_B_Mem64),
      .Data_Output_A_Mem2 (Data_Output_A_Mem65),
      .Data_Output_B_Mem2 (Data_Output_B_Mem65),
      .Data_Output_A_Mem3 (Data_Output_A_Mem66),
      .Data_Output_B_Mem3 (Data_Output_B_Mem66),
      .Data_Output_A_Mem4 (Data_Output_A_Mem67),
      .Data_Output_B_Mem4 (Data_Output_B_Mem67),
      .Data_Output_A_Mem5 (Data_Output_A_Mem68),
      .Data_Output_B_Mem5 (Data_Output_B_Mem68),
      .Data_Output_A_Mem6 (Data_Output_A_Mem69),
      .Data_Output_B_Mem6 (Data_Output_B_Mem69),
      .Data_Output_A_Mem7 (Data_Output_A_Mem70),
      .Data_Output_B_Mem7 (Data_Output_B_Mem70)
	  );
	
mem_unit #( .DATA_WIDTH(DATA_WIDTH),.IFM_SIZE(IFM_SIZE))
M11(  .clk(clk),
      .Data_Input_A_Mem1 (data_in_from_previous1),
      .Data_Input_B_Mem1 ('b0),
      .Data_Input_A_Mem2 (data_in_from_previous2),
      .Data_Input_B_Mem2 ('b0),
      .Data_Input_A_Mem3 (data_in_from_previous3),
      .Data_Input_B_Mem3 ('b0),
      .Data_Input_A_Mem4 (data_in_from_previous4),
      .Data_Input_B_Mem4 ('b0),
      .Data_Input_A_Mem5 (data_in_from_previous5),
      .Data_Input_B_Mem5 ('b0),
      .Data_Input_A_Mem6 (data_in_from_previous6),
      .Data_Input_B_Mem6 ('b0),
      .Data_Input_A_Mem7 (data_in_from_previous7),
      .Data_Input_B_Mem7 ('b0),
	
      .Address_A ( ifm_address_write_previous_dMuxOut11 | ifm_address_read_A_next_dMuxOut12 ),
      .Address_B ( ifm_address_read_previous_dMuxOut11  | ifm_address_read_B_next_dMuxOut12 ),  
	
      .Enable_Write_A_Mem (ifm_enable_write_previous_dMuxOut11),
      .Enable_Read_A_Mem  (ifm_enable_read_A_next_dMuxOut12),
      .Enable_Write_B_Mem (1'b0),
      .Enable_Read_B_Mem  (ifm_enable_read_previous_dMuxOut11 | ifm_enable_read_B_next_dMuxOut12),
	  
      .Data_Output_A_Mem1 (Data_Output_A_Mem71),
      .Data_Output_B_Mem1 (Data_Output_B_Mem71),
      .Data_Output_A_Mem2 (Data_Output_A_Mem72),
      .Data_Output_B_Mem2 (Data_Output_B_Mem72),
      .Data_Output_A_Mem3 (Data_Output_A_Mem73),
      .Data_Output_B_Mem3 (Data_Output_B_Mem73),
      .Data_Output_A_Mem4 (Data_Output_A_Mem74),
      .Data_Output_B_Mem4 (Data_Output_B_Mem74),
      .Data_Output_A_Mem5 (Data_Output_A_Mem75),
      .Data_Output_B_Mem5 (Data_Output_B_Mem75),
      .Data_Output_A_Mem6 (Data_Output_A_Mem76),
      .Data_Output_B_Mem6 (Data_Output_B_Mem76),
      .Data_Output_A_Mem7 (Data_Output_A_Mem77),
      .Data_Output_B_Mem7 (Data_Output_B_Mem77)
	  );
	
mem_unit #( .DATA_WIDTH(DATA_WIDTH),.IFM_SIZE(IFM_SIZE))
M12(  .clk(clk),
      .Data_Input_A_Mem1 (data_in_from_previous1),
      .Data_Input_B_Mem1 ('b0),
      .Data_Input_A_Mem2 (data_in_from_previous2),
      .Data_Input_B_Mem2 ('b0),
      .Data_Input_A_Mem3 (data_in_from_previous3),
      .Data_Input_B_Mem3 ('b0),
      .Data_Input_A_Mem4 (data_in_from_previous4),
      .Data_Input_B_Mem4 ('b0),
      .Data_Input_A_Mem5 (data_in_from_previous5),
      .Data_Input_B_Mem5 ('b0),
      .Data_Input_A_Mem6 (data_in_from_previous6),
      .Data_Input_B_Mem6 ('b0),
      .Data_Input_A_Mem7 (data_in_from_previous7),
      .Data_Input_B_Mem7 ('b0),
	
      .Address_A ( ifm_address_write_previous_dMuxOut12 | ifm_address_read_A_next_dMuxOut13 ),
      .Address_B ( ifm_address_read_previous_dMuxOut12  | ifm_address_read_B_next_dMuxOut13 ),  
	
      .Enable_Write_A_Mem (ifm_enable_write_previous_dMuxOut12),
      .Enable_Read_A_Mem  (ifm_enable_read_A_next_dMuxOut13),
      .Enable_Write_B_Mem (1'b0),
      .Enable_Read_B_Mem  (ifm_enable_read_previous_dMuxOut12 | ifm_enable_read_B_next_dMuxOut13),
	  
      .Data_Output_A_Mem1 (Data_Output_A_Mem78),
      .Data_Output_B_Mem1 (Data_Output_B_Mem78),
      .Data_Output_A_Mem2 (Data_Output_A_Mem79),
      .Data_Output_B_Mem2 (Data_Output_B_Mem79),
      .Data_Output_A_Mem3 (Data_Output_A_Mem80),
      .Data_Output_B_Mem3 (Data_Output_B_Mem80),
      .Data_Output_A_Mem4 (Data_Output_A_Mem81),
      .Data_Output_B_Mem4 (Data_Output_B_Mem81),
      .Data_Output_A_Mem5 (Data_Output_A_Mem82),
      .Data_Output_B_Mem5 (Data_Output_B_Mem82),
      .Data_Output_A_Mem6 (Data_Output_A_Mem83),
      .Data_Output_B_Mem6 (Data_Output_B_Mem83),
      .Data_Output_A_Mem7 (Data_Output_A_Mem84),
      .Data_Output_B_Mem7 (Data_Output_B_Mem84)
	  );
	
mem_unit #( .DATA_WIDTH(DATA_WIDTH),.IFM_SIZE(IFM_SIZE))
M13(  .clk(clk),
      .Data_Input_A_Mem1 (data_in_from_previous1),
      .Data_Input_B_Mem1 ('b0),
      .Data_Input_A_Mem2 (data_in_from_previous2),
      .Data_Input_B_Mem2 ('b0),
      .Data_Input_A_Mem3 (data_in_from_previous3),
      .Data_Input_B_Mem3 ('b0),
      .Data_Input_A_Mem4 (data_in_from_previous4),
      .Data_Input_B_Mem4 ('b0),
      .Data_Input_A_Mem5 (data_in_from_previous5),
      .Data_Input_B_Mem5 ('b0),
      .Data_Input_A_Mem6 (data_in_from_previous6),
      .Data_Input_B_Mem6 ('b0),
      .Data_Input_A_Mem7 (data_in_from_previous7),
      .Data_Input_B_Mem7 ('b0),
	
      .Address_A ( ifm_address_write_previous_dMuxOut13 | ifm_address_read_A_next_dMuxOut14 ),
      .Address_B ( ifm_address_read_previous_dMuxOut13  | ifm_address_read_B_next_dMuxOut14 ),  
	
      .Enable_Write_A_Mem (ifm_enable_write_previous_dMuxOut13),
      .Enable_Read_A_Mem  (ifm_enable_read_A_next_dMuxOut14),
      .Enable_Write_B_Mem (1'b0),
      .Enable_Read_B_Mem  (ifm_enable_read_previous_dMuxOut13 | ifm_enable_read_B_next_dMuxOut14),
	  
      .Data_Output_A_Mem1 (Data_Output_A_Mem85),
      .Data_Output_B_Mem1 (Data_Output_B_Mem85),
      .Data_Output_A_Mem2 (Data_Output_A_Mem86),
      .Data_Output_B_Mem2 (Data_Output_B_Mem86),
      .Data_Output_A_Mem3 (Data_Output_A_Mem87),
      .Data_Output_B_Mem3 (Data_Output_B_Mem87),
      .Data_Output_A_Mem4 (Data_Output_A_Mem88),
      .Data_Output_B_Mem4 (Data_Output_B_Mem88),
      .Data_Output_A_Mem5 (Data_Output_A_Mem89),
      .Data_Output_B_Mem5 (Data_Output_B_Mem89),
      .Data_Output_A_Mem6 (Data_Output_A_Mem90),
      .Data_Output_B_Mem6 (Data_Output_B_Mem90),
      .Data_Output_A_Mem7 (Data_Output_A_Mem91),
      .Data_Output_B_Mem7 (Data_Output_B_Mem91)
	  );
	
mem_unit #( .DATA_WIDTH(DATA_WIDTH),.IFM_SIZE(IFM_SIZE))
M14(  .clk(clk),
      .Data_Input_A_Mem1 (data_in_from_previous1),
      .Data_Input_B_Mem1 ('b0),
      .Data_Input_A_Mem2 (data_in_from_previous2),
      .Data_Input_B_Mem2 ('b0),
      .Data_Input_A_Mem3 (data_in_from_previous3),
      .Data_Input_B_Mem3 ('b0),
      .Data_Input_A_Mem4 (data_in_from_previous4),
      .Data_Input_B_Mem4 ('b0),
      .Data_Input_A_Mem5 (data_in_from_previous5),
      .Data_Input_B_Mem5 ('b0),
      .Data_Input_A_Mem6 (data_in_from_previous6),
      .Data_Input_B_Mem6 ('b0),
      .Data_Input_A_Mem7 (data_in_from_previous7),
      .Data_Input_B_Mem7 ('b0),
	
      .Address_A ( ifm_address_write_previous_dMuxOut14 | ifm_address_read_A_next_dMuxOut15 ),
      .Address_B ( ifm_address_read_previous_dMuxOut14  | ifm_address_read_B_next_dMuxOut15 ),  
	
      .Enable_Write_A_Mem (ifm_enable_write_previous_dMuxOut14),
      .Enable_Read_A_Mem  (ifm_enable_read_A_next_dMuxOut15),
      .Enable_Write_B_Mem (1'b0),
      .Enable_Read_B_Mem  (ifm_enable_read_previous_dMuxOut14 | ifm_enable_read_B_next_dMuxOut15),
	  
      .Data_Output_A_Mem1 (Data_Output_A_Mem92),
      .Data_Output_B_Mem1 (Data_Output_B_Mem92),
      .Data_Output_A_Mem2 (Data_Output_A_Mem93),
      .Data_Output_B_Mem2 (Data_Output_B_Mem93),
      .Data_Output_A_Mem3 (Data_Output_A_Mem94),
      .Data_Output_B_Mem3 (Data_Output_B_Mem94),
      .Data_Output_A_Mem4 (Data_Output_A_Mem95),
      .Data_Output_B_Mem4 (Data_Output_B_Mem95),
      .Data_Output_A_Mem5 (Data_Output_A_Mem96),
      .Data_Output_B_Mem5 (Data_Output_B_Mem96),
      .Data_Output_A_Mem6 (Data_Output_A_Mem97),
      .Data_Output_B_Mem6 (Data_Output_B_Mem97),
      .Data_Output_A_Mem7 (Data_Output_A_Mem98),
      .Data_Output_B_Mem7 (Data_Output_B_Mem98)
	  );
	
mem_unit #( .DATA_WIDTH(DATA_WIDTH),.IFM_SIZE(IFM_SIZE))
M15(  .clk(clk),
      .Data_Input_A_Mem1 (data_in_from_previous1),
      .Data_Input_B_Mem1 ('b0),
      .Data_Input_A_Mem2 (data_in_from_previous2),
      .Data_Input_B_Mem2 ('b0),
      .Data_Input_A_Mem3 (data_in_from_previous3),
      .Data_Input_B_Mem3 ('b0),
      .Data_Input_A_Mem4 (data_in_from_previous4),
      .Data_Input_B_Mem4 ('b0),
      .Data_Input_A_Mem5 (data_in_from_previous5),
      .Data_Input_B_Mem5 ('b0),
      .Data_Input_A_Mem6 (data_in_from_previous6),
      .Data_Input_B_Mem6 ('b0),
      .Data_Input_A_Mem7 (data_in_from_previous7),
      .Data_Input_B_Mem7 ('b0),
	
      .Address_A ( ifm_address_write_previous_dMuxOut15 | ifm_address_read_A_next_dMuxOut16 ),
      .Address_B ( ifm_address_read_previous_dMuxOut15  | ifm_address_read_B_next_dMuxOut16 ),  
	
      .Enable_Write_A_Mem (ifm_enable_write_previous_dMuxOut15),
      .Enable_Read_A_Mem  (ifm_enable_read_A_next_dMuxOut16),
      .Enable_Write_B_Mem (1'b0),
      .Enable_Read_B_Mem  (ifm_enable_read_previous_dMuxOut15 | ifm_enable_read_B_next_dMuxOut16),
	  
      .Data_Output_A_Mem1 (Data_Output_A_Mem99),
      .Data_Output_B_Mem1 (Data_Output_B_Mem99),
      .Data_Output_A_Mem2 (Data_Output_A_Mem100),
      .Data_Output_B_Mem2 (Data_Output_B_Mem100),
      .Data_Output_A_Mem3 (Data_Output_A_Mem101),
      .Data_Output_B_Mem3 (Data_Output_B_Mem101),
      .Data_Output_A_Mem4 (Data_Output_A_Mem102),
      .Data_Output_B_Mem4 (Data_Output_B_Mem102),
      .Data_Output_A_Mem5 (Data_Output_A_Mem103),
      .Data_Output_B_Mem5 (Data_Output_B_Mem103),
      .Data_Output_A_Mem6 (Data_Output_A_Mem104),
      .Data_Output_B_Mem6 (Data_Output_B_Mem104),
      .Data_Output_A_Mem7 (Data_Output_A_Mem105),
      .Data_Output_B_Mem7 (Data_Output_B_Mem105)
	  );
	
mem_unit #( .DATA_WIDTH(DATA_WIDTH),.IFM_SIZE(IFM_SIZE))
M16(  .clk(clk),
      .Data_Input_A_Mem1 (data_in_from_previous1),
      .Data_Input_B_Mem1 ('b0),
      .Data_Input_A_Mem2 (data_in_from_previous2),
      .Data_Input_B_Mem2 ('b0),
      .Data_Input_A_Mem3 (data_in_from_previous3),
      .Data_Input_B_Mem3 ('b0),
      .Data_Input_A_Mem4 (data_in_from_previous4),
      .Data_Input_B_Mem4 ('b0),
      .Data_Input_A_Mem5 (data_in_from_previous5),
      .Data_Input_B_Mem5 ('b0),
      .Data_Input_A_Mem6 (data_in_from_previous6),
      .Data_Input_B_Mem6 ('b0),
      .Data_Input_A_Mem7 (data_in_from_previous7),
      .Data_Input_B_Mem7 ('b0),
	
      .Address_A ( ifm_address_write_previous_dMuxOut16 | ifm_address_read_A_next_dMuxOut17 ),
      .Address_B ( ifm_address_read_previous_dMuxOut16  | ifm_address_read_B_next_dMuxOut17 ),  
	
      .Enable_Write_A_Mem (ifm_enable_write_previous_dMuxOut16),
      .Enable_Read_A_Mem  (ifm_enable_read_A_next_dMuxOut17),
      .Enable_Write_B_Mem (1'b0),
      .Enable_Read_B_Mem  (ifm_enable_read_previous_dMuxOut16 | ifm_enable_read_B_next_dMuxOut17),
	  
      .Data_Output_A_Mem1 (Data_Output_A_Mem106),
      .Data_Output_B_Mem1 (Data_Output_B_Mem106),
      .Data_Output_A_Mem2 (Data_Output_A_Mem107),
      .Data_Output_B_Mem2 (Data_Output_B_Mem107),
      .Data_Output_A_Mem3 (Data_Output_A_Mem108),
      .Data_Output_B_Mem3 (Data_Output_B_Mem108),
      .Data_Output_A_Mem4 (Data_Output_A_Mem109),
      .Data_Output_B_Mem4 (Data_Output_B_Mem109),
      .Data_Output_A_Mem5 (Data_Output_A_Mem110),
      .Data_Output_B_Mem5 (Data_Output_B_Mem110),
      .Data_Output_A_Mem6 (Data_Output_A_Mem111),
      .Data_Output_B_Mem6 (Data_Output_B_Mem111),
      .Data_Output_A_Mem7 (Data_Output_A_Mem112),
      .Data_Output_B_Mem7 (Data_Output_B_Mem112)
	  );
	
mem_unit #( .DATA_WIDTH(DATA_WIDTH),.IFM_SIZE(IFM_SIZE))
M17(  .clk(clk),
      .Data_Input_A_Mem1 (data_in_from_previous1),
      .Data_Input_B_Mem1 ('b0),
      .Data_Input_A_Mem2 (data_in_from_previous2),
      .Data_Input_B_Mem2 ('b0),
      .Data_Input_A_Mem3 (data_in_from_previous3),
      .Data_Input_B_Mem3 ('b0),
      .Data_Input_A_Mem4 (data_in_from_previous4),
      .Data_Input_B_Mem4 ('b0),
      .Data_Input_A_Mem5 (data_in_from_previous5),
      .Data_Input_B_Mem5 ('b0),
      .Data_Input_A_Mem6 (data_in_from_previous6),
      .Data_Input_B_Mem6 ('b0),
      .Data_Input_A_Mem7 (data_in_from_previous7),
      .Data_Input_B_Mem7 ('b0),
	
      .Address_A ( ifm_address_write_previous_dMuxOut17 | ifm_address_read_A_next_dMuxOut18 ),
      .Address_B ( ifm_address_read_previous_dMuxOut17  | ifm_address_read_B_next_dMuxOut18 ),  
	
      .Enable_Write_A_Mem (ifm_enable_write_previous_dMuxOut17),
      .Enable_Read_A_Mem  (ifm_enable_read_A_next_dMuxOut18),
      .Enable_Write_B_Mem (1'b0),
      .Enable_Read_B_Mem  (ifm_enable_read_previous_dMuxOut17 | ifm_enable_read_B_next_dMuxOut18),
	  
      .Data_Output_A_Mem1 (Data_Output_A_Mem113),
      .Data_Output_B_Mem1 (Data_Output_B_Mem113),
      .Data_Output_A_Mem2 (Data_Output_A_Mem114),
      .Data_Output_B_Mem2 (Data_Output_B_Mem114),
      .Data_Output_A_Mem3 (Data_Output_A_Mem115),
      .Data_Output_B_Mem3 (Data_Output_B_Mem115),
      .Data_Output_A_Mem4 (Data_Output_A_Mem116),
      .Data_Output_B_Mem4 (Data_Output_B_Mem116),
      .Data_Output_A_Mem5 (Data_Output_A_Mem117),
      .Data_Output_B_Mem5 (Data_Output_B_Mem117),
      .Data_Output_A_Mem6 (Data_Output_A_Mem118),
      .Data_Output_B_Mem6 (Data_Output_B_Mem118),
      .Data_Output_A_Mem7 (Data_Output_A_Mem119),
      .Data_Output_B_Mem7 (Data_Output_B_Mem119)
	  );
	
mem_unit #( .DATA_WIDTH(DATA_WIDTH),.IFM_SIZE(IFM_SIZE))
M18(  .clk(clk),
      .Data_Input_A_Mem1 (data_in_from_previous1),
      .Data_Input_B_Mem1 ('b0),
      .Data_Input_A_Mem2 (data_in_from_previous2),
      .Data_Input_B_Mem2 ('b0),
      .Data_Input_A_Mem3 (data_in_from_previous3),
      .Data_Input_B_Mem3 ('b0),
      .Data_Input_A_Mem4 (data_in_from_previous4),
      .Data_Input_B_Mem4 ('b0),
      .Data_Input_A_Mem5 (data_in_from_previous5),
      .Data_Input_B_Mem5 ('b0),
      .Data_Input_A_Mem6 (data_in_from_previous6),
      .Data_Input_B_Mem6 ('b0),
      .Data_Input_A_Mem7 (data_in_from_previous7),
      .Data_Input_B_Mem7 ('b0),
	
      .Address_A ( ifm_address_write_previous_dMuxOut18 | ifm_address_read_A_next_dMuxOut19 ),
      .Address_B ( ifm_address_read_previous_dMuxOut18  | ifm_address_read_B_next_dMuxOut19 ),  
	
      .Enable_Write_A_Mem (ifm_enable_write_previous_dMuxOut18),
      .Enable_Read_A_Mem  (ifm_enable_read_A_next_dMuxOut19),
      .Enable_Write_B_Mem (1'b0),
      .Enable_Read_B_Mem  (ifm_enable_read_previous_dMuxOut18 | ifm_enable_read_B_next_dMuxOut19),
	  
      .Data_Output_A_Mem1 (Data_Output_A_Mem120),
      .Data_Output_B_Mem1 (Data_Output_B_Mem120),
      .Data_Output_A_Mem2 (Data_Output_A_Mem121),
      .Data_Output_B_Mem2 (Data_Output_B_Mem121),
      .Data_Output_A_Mem3 (Data_Output_A_Mem122),
      .Data_Output_B_Mem3 (Data_Output_B_Mem122),
      .Data_Output_A_Mem4 (Data_Output_A_Mem123),
      .Data_Output_B_Mem4 (Data_Output_B_Mem123),
      .Data_Output_A_Mem5 (Data_Output_A_Mem124),
      .Data_Output_B_Mem5 (Data_Output_B_Mem124),
      .Data_Output_A_Mem6 (Data_Output_A_Mem125),
      .Data_Output_B_Mem6 (Data_Output_B_Mem125),
      .Data_Output_A_Mem7 (Data_Output_A_Mem126),
      .Data_Output_B_Mem7 (Data_Output_B_Mem126)
	  );
	
mem_unit #( .DATA_WIDTH(DATA_WIDTH),.IFM_SIZE(IFM_SIZE))
M19(  .clk(clk),
      .Data_Input_A_Mem1 (data_in_from_previous1),
      .Data_Input_B_Mem1 ('b0),
      .Data_Input_A_Mem2 (data_in_from_previous2),
      .Data_Input_B_Mem2 ('b0),
      .Data_Input_A_Mem3 (data_in_from_previous3),
      .Data_Input_B_Mem3 ('b0),
      .Data_Input_A_Mem4 (data_in_from_previous4),
      .Data_Input_B_Mem4 ('b0),
      .Data_Input_A_Mem5 (data_in_from_previous5),
      .Data_Input_B_Mem5 ('b0),
      .Data_Input_A_Mem6 (data_in_from_previous6),
      .Data_Input_B_Mem6 ('b0),
      .Data_Input_A_Mem7 (data_in_from_previous7),
      .Data_Input_B_Mem7 ('b0),
	
      .Address_A ( ifm_address_write_previous_dMuxOut19 | ifm_address_read_A_next_dMuxOut20 ),
      .Address_B ( ifm_address_read_previous_dMuxOut19  | ifm_address_read_B_next_dMuxOut20 ),  
	
      .Enable_Write_A_Mem (ifm_enable_write_previous_dMuxOut19),
      .Enable_Read_A_Mem  (ifm_enable_read_A_next_dMuxOut20),
      .Enable_Write_B_Mem (1'b0),
      .Enable_Read_B_Mem  (ifm_enable_read_previous_dMuxOut19 | ifm_enable_read_B_next_dMuxOut20),
	  
      .Data_Output_A_Mem1 (Data_Output_A_Mem127),
      .Data_Output_B_Mem1 (Data_Output_B_Mem127),
      .Data_Output_A_Mem2 (Data_Output_A_Mem128),
      .Data_Output_B_Mem2 (Data_Output_B_Mem128),
      .Data_Output_A_Mem3 (Data_Output_A_Mem129),
      .Data_Output_B_Mem3 (Data_Output_B_Mem129),
      .Data_Output_A_Mem4 (Data_Output_A_Mem130),
      .Data_Output_B_Mem4 (Data_Output_B_Mem130),
      .Data_Output_A_Mem5 (Data_Output_A_Mem131),
      .Data_Output_B_Mem5 (Data_Output_B_Mem131),
      .Data_Output_A_Mem6 (Data_Output_A_Mem132),
      .Data_Output_B_Mem6 (Data_Output_B_Mem132),
      .Data_Output_A_Mem7 (Data_Output_A_Mem133),
      .Data_Output_B_Mem7 (Data_Output_B_Mem133)
	  );
	
mem_unit #( .DATA_WIDTH(DATA_WIDTH),.IFM_SIZE(IFM_SIZE))
M20(  .clk(clk),
      .Data_Input_A_Mem1 (data_in_from_previous1),
      .Data_Input_B_Mem1 ('b0),
      .Data_Input_A_Mem2 (data_in_from_previous2),
      .Data_Input_B_Mem2 ('b0),
      .Data_Input_A_Mem3 (data_in_from_previous3),
      .Data_Input_B_Mem3 ('b0),
      .Data_Input_A_Mem4 (data_in_from_previous4),
      .Data_Input_B_Mem4 ('b0),
      .Data_Input_A_Mem5 (data_in_from_previous5),
      .Data_Input_B_Mem5 ('b0),
      .Data_Input_A_Mem6 (data_in_from_previous6),
      .Data_Input_B_Mem6 ('b0),
      .Data_Input_A_Mem7 (data_in_from_previous7),
      .Data_Input_B_Mem7 ('b0),
	
      .Address_A ( ifm_address_write_previous_dMuxOut20 | ifm_address_read_A_next_dMuxOut21 ),
      .Address_B ( ifm_address_read_previous_dMuxOut20  | ifm_address_read_B_next_dMuxOut21 ),  
	
      .Enable_Write_A_Mem (ifm_enable_write_previous_dMuxOut20),
      .Enable_Read_A_Mem  (ifm_enable_read_A_next_dMuxOut21),
      .Enable_Write_B_Mem (1'b0),
      .Enable_Read_B_Mem  (ifm_enable_read_previous_dMuxOut20 | ifm_enable_read_B_next_dMuxOut21),
	  
      .Data_Output_A_Mem1 (Data_Output_A_Mem134),
      .Data_Output_B_Mem1 (Data_Output_B_Mem134),
      .Data_Output_A_Mem2 (Data_Output_A_Mem135),
      .Data_Output_B_Mem2 (Data_Output_B_Mem135),
      .Data_Output_A_Mem3 (Data_Output_A_Mem136),
      .Data_Output_B_Mem3 (Data_Output_B_Mem136),
      .Data_Output_A_Mem4 (Data_Output_A_Mem137),
      .Data_Output_B_Mem4 (Data_Output_B_Mem137),
      .Data_Output_A_Mem5 (Data_Output_A_Mem138),
      .Data_Output_B_Mem5 (Data_Output_B_Mem138),
      .Data_Output_A_Mem6 (Data_Output_A_Mem139),
      .Data_Output_B_Mem6 (Data_Output_B_Mem139),
      .Data_Output_A_Mem7 (Data_Output_A_Mem140),
      .Data_Output_B_Mem7 (Data_Output_B_Mem140)
	  );
	
mem_unit #( .DATA_WIDTH(DATA_WIDTH),.IFM_SIZE(IFM_SIZE))
M21(  .clk(clk),
      .Data_Input_A_Mem1 (data_in_from_previous1),
      .Data_Input_B_Mem1 ('b0),
      .Data_Input_A_Mem2 (data_in_from_previous2),
      .Data_Input_B_Mem2 ('b0),
      .Data_Input_A_Mem3 (data_in_from_previous3),
      .Data_Input_B_Mem3 ('b0),
      .Data_Input_A_Mem4 (data_in_from_previous4),
      .Data_Input_B_Mem4 ('b0),
      .Data_Input_A_Mem5 (data_in_from_previous5),
      .Data_Input_B_Mem5 ('b0),
      .Data_Input_A_Mem6 (data_in_from_previous6),
      .Data_Input_B_Mem6 ('b0),
      .Data_Input_A_Mem7 (data_in_from_previous7),
      .Data_Input_B_Mem7 ('b0),
	
      .Address_A ( ifm_address_write_previous_dMuxOut21 | ifm_address_read_A_next_dMuxOut22 ),
      .Address_B ( ifm_address_read_previous_dMuxOut21  | ifm_address_read_B_next_dMuxOut22 ),  
	
      .Enable_Write_A_Mem (ifm_enable_write_previous_dMuxOut21),
      .Enable_Read_A_Mem  (ifm_enable_read_A_next_dMuxOut22),
      .Enable_Write_B_Mem (1'b0),
      .Enable_Read_B_Mem  (ifm_enable_read_previous_dMuxOut21 | ifm_enable_read_B_next_dMuxOut22),
	  
      .Data_Output_A_Mem1 (Data_Output_A_Mem141),
      .Data_Output_B_Mem1 (Data_Output_B_Mem141),
      .Data_Output_A_Mem2 (Data_Output_A_Mem142),
      .Data_Output_B_Mem2 (Data_Output_B_Mem142),
      .Data_Output_A_Mem3 (Data_Output_A_Mem143),
      .Data_Output_B_Mem3 (Data_Output_B_Mem143),
      .Data_Output_A_Mem4 (Data_Output_A_Mem144),
      .Data_Output_B_Mem4 (Data_Output_B_Mem144),
      .Data_Output_A_Mem5 (Data_Output_A_Mem145),
      .Data_Output_B_Mem5 (Data_Output_B_Mem145),
      .Data_Output_A_Mem6 (Data_Output_A_Mem146),
      .Data_Output_B_Mem6 (Data_Output_B_Mem146),
      .Data_Output_A_Mem7 (Data_Output_A_Mem147),
      .Data_Output_B_Mem7 (Data_Output_B_Mem147)
	  );
	
mem_unit #( .DATA_WIDTH(DATA_WIDTH),.IFM_SIZE(IFM_SIZE))
M22(  .clk(clk),
      .Data_Input_A_Mem1 (data_in_from_previous1),
      .Data_Input_B_Mem1 ('b0),
      .Data_Input_A_Mem2 (data_in_from_previous2),
      .Data_Input_B_Mem2 ('b0),
      .Data_Input_A_Mem3 (data_in_from_previous3),
      .Data_Input_B_Mem3 ('b0),
      .Data_Input_A_Mem4 (data_in_from_previous4),
      .Data_Input_B_Mem4 ('b0),
      .Data_Input_A_Mem5 (data_in_from_previous5),
      .Data_Input_B_Mem5 ('b0),
      .Data_Input_A_Mem6 (data_in_from_previous6),
      .Data_Input_B_Mem6 ('b0),
      .Data_Input_A_Mem7 (data_in_from_previous7),
      .Data_Input_B_Mem7 ('b0),
	
      .Address_A ( ifm_address_write_previous_dMuxOut22 | ifm_address_read_A_next_dMuxOut23 ),
      .Address_B ( ifm_address_read_previous_dMuxOut22  | ifm_address_read_B_next_dMuxOut23 ),  
	
      .Enable_Write_A_Mem (ifm_enable_write_previous_dMuxOut22),
      .Enable_Read_A_Mem  (ifm_enable_read_A_next_dMuxOut23),
      .Enable_Write_B_Mem (1'b0),
      .Enable_Read_B_Mem  (ifm_enable_read_previous_dMuxOut22 | ifm_enable_read_B_next_dMuxOut23),
	  
      .Data_Output_A_Mem1 (Data_Output_A_Mem148),
      .Data_Output_B_Mem1 (Data_Output_B_Mem148),
      .Data_Output_A_Mem2 (Data_Output_A_Mem149),
      .Data_Output_B_Mem2 (Data_Output_B_Mem149),
      .Data_Output_A_Mem3 (Data_Output_A_Mem150),
      .Data_Output_B_Mem3 (Data_Output_B_Mem150),
      .Data_Output_A_Mem4 (Data_Output_A_Mem151),
      .Data_Output_B_Mem4 (Data_Output_B_Mem151),
      .Data_Output_A_Mem5 (Data_Output_A_Mem152),
      .Data_Output_B_Mem5 (Data_Output_B_Mem152),
      .Data_Output_A_Mem6 (Data_Output_A_Mem153),
      .Data_Output_B_Mem6 (Data_Output_B_Mem153),
      .Data_Output_A_Mem7 (Data_Output_A_Mem154),
      .Data_Output_B_Mem7 (Data_Output_B_Mem154)
	  );
	
mem_unit #( .DATA_WIDTH(DATA_WIDTH),.IFM_SIZE(IFM_SIZE))
M23(  .clk(clk),
      .Data_Input_A_Mem1 (data_in_from_previous1),
      .Data_Input_B_Mem1 ('b0),
      .Data_Input_A_Mem2 (data_in_from_previous2),
      .Data_Input_B_Mem2 ('b0),
      .Data_Input_A_Mem3 (data_in_from_previous3),
      .Data_Input_B_Mem3 ('b0),
      .Data_Input_A_Mem4 (data_in_from_previous4),
      .Data_Input_B_Mem4 ('b0),
      .Data_Input_A_Mem5 (data_in_from_previous5),
      .Data_Input_B_Mem5 ('b0),
      .Data_Input_A_Mem6 (data_in_from_previous6),
      .Data_Input_B_Mem6 ('b0),
      .Data_Input_A_Mem7 (data_in_from_previous7),
      .Data_Input_B_Mem7 ('b0),
	
      .Address_A ( ifm_address_write_previous_dMuxOut23 | ifm_address_read_A_next_dMuxOut24 ),
      .Address_B ( ifm_address_read_previous_dMuxOut23  | ifm_address_read_B_next_dMuxOut24 ),  
	
      .Enable_Write_A_Mem (ifm_enable_write_previous_dMuxOut23),
      .Enable_Read_A_Mem  (ifm_enable_read_A_next_dMuxOut24),
      .Enable_Write_B_Mem (1'b0),
      .Enable_Read_B_Mem  (ifm_enable_read_previous_dMuxOut23 | ifm_enable_read_B_next_dMuxOut24),
	  
      .Data_Output_A_Mem1 (Data_Output_A_Mem155),
      .Data_Output_B_Mem1 (Data_Output_B_Mem155),
      .Data_Output_A_Mem2 (Data_Output_A_Mem156),
      .Data_Output_B_Mem2 (Data_Output_B_Mem156),
      .Data_Output_A_Mem3 (Data_Output_A_Mem157),
      .Data_Output_B_Mem3 (Data_Output_B_Mem157),
      .Data_Output_A_Mem4 (Data_Output_A_Mem158),
      .Data_Output_B_Mem4 (Data_Output_B_Mem158),
      .Data_Output_A_Mem5 (Data_Output_A_Mem159),
      .Data_Output_B_Mem5 (Data_Output_B_Mem159),
      .Data_Output_A_Mem6 (Data_Output_A_Mem160),
      .Data_Output_B_Mem6 (Data_Output_B_Mem160),
      .Data_Output_A_Mem7 (Data_Output_A_Mem161),
      .Data_Output_B_Mem7 (Data_Output_B_Mem161)
	  );
	
mem_unit #( .DATA_WIDTH(DATA_WIDTH),.IFM_SIZE(IFM_SIZE))
M24(  .clk(clk),
      .Data_Input_A_Mem1 (data_in_from_previous1),
      .Data_Input_B_Mem1 ('b0),
      .Data_Input_A_Mem2 (data_in_from_previous2),
      .Data_Input_B_Mem2 ('b0),
      .Data_Input_A_Mem3 (data_in_from_previous3),
      .Data_Input_B_Mem3 ('b0),
      .Data_Input_A_Mem4 (data_in_from_previous4),
      .Data_Input_B_Mem4 ('b0),
      .Data_Input_A_Mem5 (data_in_from_previous5),
      .Data_Input_B_Mem5 ('b0),
      .Data_Input_A_Mem6 (data_in_from_previous6),
      .Data_Input_B_Mem6 ('b0),
      .Data_Input_A_Mem7 (data_in_from_previous7),
      .Data_Input_B_Mem7 ('b0),
	
      .Address_A ( ifm_address_write_previous_dMuxOut24 | ifm_address_read_A_next_dMuxOut25 ),
      .Address_B ( ifm_address_read_previous_dMuxOut24  | ifm_address_read_B_next_dMuxOut25 ),  
	
      .Enable_Write_A_Mem (ifm_enable_write_previous_dMuxOut24),
      .Enable_Read_A_Mem  (ifm_enable_read_A_next_dMuxOut25),
      .Enable_Write_B_Mem (1'b0),
      .Enable_Read_B_Mem  (ifm_enable_read_previous_dMuxOut24 | ifm_enable_read_B_next_dMuxOut25),
	  
      .Data_Output_A_Mem1 (Data_Output_A_Mem162),
      .Data_Output_B_Mem1 (Data_Output_B_Mem162),
      .Data_Output_A_Mem2 (Data_Output_A_Mem163),
      .Data_Output_B_Mem2 (Data_Output_B_Mem163),
      .Data_Output_A_Mem3 (Data_Output_A_Mem164),
      .Data_Output_B_Mem3 (Data_Output_B_Mem164),
      .Data_Output_A_Mem4 (Data_Output_A_Mem165),
      .Data_Output_B_Mem4 (Data_Output_B_Mem165),
      .Data_Output_A_Mem5 (Data_Output_A_Mem166),
      .Data_Output_B_Mem5 (Data_Output_B_Mem166),
      .Data_Output_A_Mem6 (Data_Output_A_Mem167),
      .Data_Output_B_Mem6 (Data_Output_B_Mem167),
      .Data_Output_A_Mem7 (Data_Output_A_Mem168),
      .Data_Output_B_Mem7 (Data_Output_B_Mem168)
	  );
	
mem_unit #( .DATA_WIDTH(DATA_WIDTH),.IFM_SIZE(IFM_SIZE))
M25(  .clk(clk),
      .Data_Input_A_Mem1 (data_in_from_previous1),
      .Data_Input_B_Mem1 ('b0),
      .Data_Input_A_Mem2 (data_in_from_previous2),
      .Data_Input_B_Mem2 ('b0),
      .Data_Input_A_Mem3 (data_in_from_previous3),
      .Data_Input_B_Mem3 ('b0),
      .Data_Input_A_Mem4 (data_in_from_previous4),
      .Data_Input_B_Mem4 ('b0),
      .Data_Input_A_Mem5 (data_in_from_previous5),
      .Data_Input_B_Mem5 ('b0),
      .Data_Input_A_Mem6 (data_in_from_previous6),
      .Data_Input_B_Mem6 ('b0),
      .Data_Input_A_Mem7 (data_in_from_previous7),
      .Data_Input_B_Mem7 ('b0),
	
      .Address_A ( ifm_address_write_previous_dMuxOut25 | ifm_address_read_A_next_dMuxOut26 ),
      .Address_B ( ifm_address_read_previous_dMuxOut25  | ifm_address_read_B_next_dMuxOut26 ),  
	
      .Enable_Write_A_Mem (ifm_enable_write_previous_dMuxOut25),
      .Enable_Read_A_Mem  (ifm_enable_read_A_next_dMuxOut26),
      .Enable_Write_B_Mem (1'b0),
      .Enable_Read_B_Mem  (ifm_enable_read_previous_dMuxOut25 | ifm_enable_read_B_next_dMuxOut26),
	  
      .Data_Output_A_Mem1 (Data_Output_A_Mem169),
      .Data_Output_B_Mem1 (Data_Output_B_Mem169),
      .Data_Output_A_Mem2 (Data_Output_A_Mem170),
      .Data_Output_B_Mem2 (Data_Output_B_Mem170),
      .Data_Output_A_Mem3 (Data_Output_A_Mem171),
      .Data_Output_B_Mem3 (Data_Output_B_Mem171),
      .Data_Output_A_Mem4 (Data_Output_A_Mem172),
      .Data_Output_B_Mem4 (Data_Output_B_Mem172),
      .Data_Output_A_Mem5 (Data_Output_A_Mem173),
      .Data_Output_B_Mem5 (Data_Output_B_Mem173),
      .Data_Output_A_Mem6 (Data_Output_A_Mem174),
      .Data_Output_B_Mem6 (Data_Output_B_Mem174),
      .Data_Output_A_Mem7 (Data_Output_A_Mem175),
      .Data_Output_B_Mem7 (Data_Output_B_Mem175)
	  );
	
mem_unit #( .DATA_WIDTH(DATA_WIDTH),.IFM_SIZE(IFM_SIZE))
M26(  .clk(clk),
      .Data_Input_A_Mem1 (data_in_from_previous1),
      .Data_Input_B_Mem1 ('b0),
      .Data_Input_A_Mem2 (data_in_from_previous2),
      .Data_Input_B_Mem2 ('b0),
      .Data_Input_A_Mem3 (data_in_from_previous3),
      .Data_Input_B_Mem3 ('b0),
      .Data_Input_A_Mem4 (data_in_from_previous4),
      .Data_Input_B_Mem4 ('b0),
      .Data_Input_A_Mem5 (data_in_from_previous5),
      .Data_Input_B_Mem5 ('b0),
      .Data_Input_A_Mem6 (data_in_from_previous6),
      .Data_Input_B_Mem6 ('b0),
      .Data_Input_A_Mem7 (data_in_from_previous7),
      .Data_Input_B_Mem7 ('b0),
	
      .Address_A ( ifm_address_write_previous_dMuxOut26 | ifm_address_read_A_next_dMuxOut27 ),
      .Address_B ( ifm_address_read_previous_dMuxOut26  | ifm_address_read_B_next_dMuxOut27 ),  
	
      .Enable_Write_A_Mem (ifm_enable_write_previous_dMuxOut26),
      .Enable_Read_A_Mem  (ifm_enable_read_A_next_dMuxOut27),
      .Enable_Write_B_Mem (1'b0),
      .Enable_Read_B_Mem  (ifm_enable_read_previous_dMuxOut26 | ifm_enable_read_B_next_dMuxOut27),
	  
      .Data_Output_A_Mem1 (Data_Output_A_Mem176),
      .Data_Output_B_Mem1 (Data_Output_B_Mem176),
      .Data_Output_A_Mem2 (Data_Output_A_Mem177),
      .Data_Output_B_Mem2 (Data_Output_B_Mem177),
      .Data_Output_A_Mem3 (Data_Output_A_Mem178),
      .Data_Output_B_Mem3 (Data_Output_B_Mem178),
      .Data_Output_A_Mem4 (Data_Output_A_Mem179),
      .Data_Output_B_Mem4 (Data_Output_B_Mem179),
      .Data_Output_A_Mem5 (Data_Output_A_Mem180),
      .Data_Output_B_Mem5 (Data_Output_B_Mem180),
      .Data_Output_A_Mem6 (Data_Output_A_Mem181),
      .Data_Output_B_Mem6 (Data_Output_B_Mem181),
      .Data_Output_A_Mem7 (Data_Output_A_Mem182),
      .Data_Output_B_Mem7 (Data_Output_B_Mem182)
	  );
	
mem_unit #( .DATA_WIDTH(DATA_WIDTH),.IFM_SIZE(IFM_SIZE))
M27(  .clk(clk),
      .Data_Input_A_Mem1 (data_in_from_previous1),
      .Data_Input_B_Mem1 ('b0),
      .Data_Input_A_Mem2 (data_in_from_previous2),
      .Data_Input_B_Mem2 ('b0),
      .Data_Input_A_Mem3 (data_in_from_previous3),
      .Data_Input_B_Mem3 ('b0),
      .Data_Input_A_Mem4 (data_in_from_previous4),
      .Data_Input_B_Mem4 ('b0),
      .Data_Input_A_Mem5 (data_in_from_previous5),
      .Data_Input_B_Mem5 ('b0),
      .Data_Input_A_Mem6 (data_in_from_previous6),
      .Data_Input_B_Mem6 ('b0),
      .Data_Input_A_Mem7 (data_in_from_previous7),
      .Data_Input_B_Mem7 ('b0),
	
      .Address_A ( ifm_address_write_previous_dMuxOut27 | ifm_address_read_A_next_dMuxOut28 ),
      .Address_B ( ifm_address_read_previous_dMuxOut27  | ifm_address_read_B_next_dMuxOut28 ),  
	
      .Enable_Write_A_Mem (ifm_enable_write_previous_dMuxOut27),
      .Enable_Read_A_Mem  (ifm_enable_read_A_next_dMuxOut28),
      .Enable_Write_B_Mem (1'b0),
      .Enable_Read_B_Mem  (ifm_enable_read_previous_dMuxOut27 | ifm_enable_read_B_next_dMuxOut28),
	  
      .Data_Output_A_Mem1 (Data_Output_A_Mem183),
      .Data_Output_B_Mem1 (Data_Output_B_Mem183),
      .Data_Output_A_Mem2 (Data_Output_A_Mem184),
      .Data_Output_B_Mem2 (Data_Output_B_Mem184),
      .Data_Output_A_Mem3 (Data_Output_A_Mem185),
      .Data_Output_B_Mem3 (Data_Output_B_Mem185),
      .Data_Output_A_Mem4 (Data_Output_A_Mem186),
      .Data_Output_B_Mem4 (Data_Output_B_Mem186),
      .Data_Output_A_Mem5 (Data_Output_A_Mem187),
      .Data_Output_B_Mem5 (Data_Output_B_Mem187),
      .Data_Output_A_Mem6 (Data_Output_A_Mem188),
      .Data_Output_B_Mem6 (Data_Output_B_Mem188),
      .Data_Output_A_Mem7 (Data_Output_A_Mem189),
      .Data_Output_B_Mem7 (Data_Output_B_Mem189)
	  );
	
mem_unit #( .DATA_WIDTH(DATA_WIDTH),.IFM_SIZE(IFM_SIZE))
M28(  .clk(clk),
      .Data_Input_A_Mem1 (data_in_from_previous1),
      .Data_Input_B_Mem1 ('b0),
      .Data_Input_A_Mem2 (data_in_from_previous2),
      .Data_Input_B_Mem2 ('b0),
      .Data_Input_A_Mem3 (data_in_from_previous3),
      .Data_Input_B_Mem3 ('b0),
      .Data_Input_A_Mem4 (data_in_from_previous4),
      .Data_Input_B_Mem4 ('b0),
      .Data_Input_A_Mem5 (data_in_from_previous5),
      .Data_Input_B_Mem5 ('b0),
      .Data_Input_A_Mem6 (data_in_from_previous6),
      .Data_Input_B_Mem6 ('b0),
      .Data_Input_A_Mem7 (data_in_from_previous7),
      .Data_Input_B_Mem7 ('b0),
	
      .Address_A ( ifm_address_write_previous_dMuxOut28 | ifm_address_read_A_next_dMuxOut29 ),
      .Address_B ( ifm_address_read_previous_dMuxOut28  | ifm_address_read_B_next_dMuxOut29 ),  
	
      .Enable_Write_A_Mem (ifm_enable_write_previous_dMuxOut28),
      .Enable_Read_A_Mem  (ifm_enable_read_A_next_dMuxOut29),
      .Enable_Write_B_Mem (1'b0),
      .Enable_Read_B_Mem  (ifm_enable_read_previous_dMuxOut28 | ifm_enable_read_B_next_dMuxOut29),
	  
      .Data_Output_A_Mem1 (Data_Output_A_Mem190),
      .Data_Output_B_Mem1 (Data_Output_B_Mem190),
      .Data_Output_A_Mem2 (Data_Output_A_Mem191),
      .Data_Output_B_Mem2 (Data_Output_B_Mem191),
      .Data_Output_A_Mem3 (Data_Output_A_Mem192),
      .Data_Output_B_Mem3 (Data_Output_B_Mem192),
      .Data_Output_A_Mem4 (Data_Output_A_Mem193),
      .Data_Output_B_Mem4 (Data_Output_B_Mem193),
      .Data_Output_A_Mem5 (Data_Output_A_Mem194),
      .Data_Output_B_Mem5 (Data_Output_B_Mem194),
      .Data_Output_A_Mem6 (Data_Output_A_Mem195),
      .Data_Output_B_Mem6 (Data_Output_B_Mem195),
      .Data_Output_A_Mem7 (Data_Output_A_Mem196),
      .Data_Output_B_Mem7 (Data_Output_B_Mem196)
	  );
	TrueDualPort_Memory #(.DATA_WIDTH(DATA_WIDTH), .MEM_SIZE(IFM_SIZE*IFM_SIZE)) 
	IFM197 (
    .clk(clk),
	
	.Data_Input_A(data_in_from_previous1),
	.Data_Input_B('b0),
	
	.Address_A ( ifm_address_write_previous_dMuxOut29 | ifm_address_read_A_next_dMuxOut1 ),
    .Address_B ( ifm_address_read_previous_dMuxOut29  | ifm_address_read_B_next_dMuxOut1 ),  
	
	.Enable_Write_A_Mem (ifm_enable_write_previous_dMuxOut29),
    .Enable_Read_A_Mem  (ifm_enable_read_A_next_dMuxOut1),
    .Enable_Write_B_Mem (1'b0),
    .Enable_Read_B_Mem  (ifm_enable_read_previous_dMuxOut29 | ifm_enable_read_B_next_dMuxOut1),
	  
	
    .Data_Output_A(Data_Output_A_Mem197),
    .Data_Output_B(Data_Output_B_Mem197)
	);
	
	TrueDualPort_Memory #(.DATA_WIDTH(DATA_WIDTH), .MEM_SIZE(IFM_SIZE*IFM_SIZE)) 
	IFM198 (
    .clk(clk),
	
	.Data_Input_A(data_in_from_previous2),
	.Data_Input_B('b0),
	
	.Address_A ( ifm_address_write_previous_dMuxOut29 | ifm_address_read_A_next_dMuxOut1 ),
    .Address_B ( ifm_address_read_previous_dMuxOut29  | ifm_address_read_B_next_dMuxOut1 ),  
	
	.Enable_Write_A_Mem (ifm_enable_write_previous_dMuxOut29),
    .Enable_Read_A_Mem  (ifm_enable_read_A_next_dMuxOut1),
    .Enable_Write_B_Mem (1'b0),
    .Enable_Read_B_Mem  (ifm_enable_read_previous_dMuxOut29 | ifm_enable_read_B_next_dMuxOut1),
	  
	
    .Data_Output_A(Data_Output_A_Mem198),
    .Data_Output_B(Data_Output_B_Mem198)
	);
	
	TrueDualPort_Memory #(.DATA_WIDTH(DATA_WIDTH), .MEM_SIZE(IFM_SIZE*IFM_SIZE)) 
	IFM199 (
    .clk(clk),
	
	.Data_Input_A(data_in_from_previous3),
	.Data_Input_B('b0),
	
	.Address_A ( ifm_address_write_previous_dMuxOut29 | ifm_address_read_A_next_dMuxOut1 ),
    .Address_B ( ifm_address_read_previous_dMuxOut29  | ifm_address_read_B_next_dMuxOut1 ),  
	
	.Enable_Write_A_Mem (ifm_enable_write_previous_dMuxOut29),
    .Enable_Read_A_Mem  (ifm_enable_read_A_next_dMuxOut1),
    .Enable_Write_B_Mem (1'b0),
    .Enable_Read_B_Mem  (ifm_enable_read_previous_dMuxOut29 | ifm_enable_read_B_next_dMuxOut1),
	  
	
    .Data_Output_A(Data_Output_A_Mem199),
    .Data_Output_B(Data_Output_B_Mem199)
	);
	
	TrueDualPort_Memory #(.DATA_WIDTH(DATA_WIDTH), .MEM_SIZE(IFM_SIZE*IFM_SIZE)) 
	IFM200 (
    .clk(clk),
	
	.Data_Input_A(data_in_from_previous4),
	.Data_Input_B('b0),
	
	.Address_A ( ifm_address_write_previous_dMuxOut29 | ifm_address_read_A_next_dMuxOut1 ),
    .Address_B ( ifm_address_read_previous_dMuxOut29  | ifm_address_read_B_next_dMuxOut1 ),  
	
	.Enable_Write_A_Mem (ifm_enable_write_previous_dMuxOut29),
    .Enable_Read_A_Mem  (ifm_enable_read_A_next_dMuxOut1),
    .Enable_Write_B_Mem (1'b0),
    .Enable_Read_B_Mem  (ifm_enable_read_previous_dMuxOut29 | ifm_enable_read_B_next_dMuxOut1),
	  
	
    .Data_Output_A(Data_Output_A_Mem200),
    .Data_Output_B(Data_Output_B_Mem200)
	);
	
endmodule